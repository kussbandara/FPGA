-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 16 2020 17:40:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SPI" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SPI
entity SPI is
port (
    ch5_B : in std_logic;
    PWM6 : out std_logic;
    ch3_A : in std_logic;
    ch0_B : in std_logic;
    PWM1 : out std_logic;
    ch4_B : in std_logic;
    RST : in std_logic;
    PWM0 : out std_logic;
    MOSI : in std_logic;
    ch7_B : in std_logic;
    PWM3 : out std_logic;
    ch2_B : in std_logic;
    SSEL : in std_logic;
    PWM2 : out std_logic;
    MISO : out std_logic;
    ch6_B : in std_logic;
    ch2_A : in std_logic;
    PWM5 : out std_logic;
    ch7_A : in std_logic;
    ch6_A : in std_logic;
    ch3_B : in std_logic;
    ch1_A : in std_logic;
    ch0_A : in std_logic;
    SCK : in std_logic;
    PWM4 : out std_logic;
    CLK : in std_logic;
    ch5_A : in std_logic;
    ch4_A : in std_logic;
    ch1_B : in std_logic;
    PWM7 : out std_logic);
end SPI;

-- Architecture of SPI
-- View name is \INTERFACE\
architecture \INTERFACE\ of SPI is

signal \N__39370\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \CLK_c\ : std_logic;
signal \PWMInstance7.un1_periodCounter12_1_0_a2_0_6_cascade_\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_0\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_1\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_2\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_3\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_4\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_5\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_6\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_7\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_8\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_9\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_10\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_11\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_12\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_13\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_14\ : std_logic;
signal \PWMInstance7.un1_periodCounter_2_cry_15\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_16\ : std_logic;
signal \PWMInstance7.periodCounter12\ : std_logic;
signal \PWMInstance7.clkCountZ0Z_0\ : std_logic;
signal \PWMInstance7.clkCountZ0Z_1\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_2\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_2\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_3\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_11\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_10\ : std_logic;
signal \PWMInstance7.un1_periodCounter12_1_0_a2_0_0\ : std_logic;
signal \PWMInstance7.un1_periodCounter12_1_0_a2_0_10\ : std_logic;
signal \PWMInstance7.un1_periodCounter12_1_0_a2_0_9\ : std_logic;
signal \PWMInstance7.un1_periodCounter12_1_0_a2_0_12_cascade_\ : std_logic;
signal \PWMInstance7.un1_periodCounter12_1_0_a2_0_14\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_4\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_5\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_8\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_9\ : std_logic;
signal \bfn_3_10_0_\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_6\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_0\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_6\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_1\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_2\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_6\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_3\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_6\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_4\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_5\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_6\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_7\ : std_logic;
signal \PWMInstance7.un1_periodCounter12_1_0_a2_0\ : std_logic;
signal \PWMInstance7.out_0_sqmuxa\ : std_logic;
signal \bfn_3_11_0_\ : std_logic;
signal \PWM7_c\ : std_logic;
signal \pwmWrite_fastZ0Z_7\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_9\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_10\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_3\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_15\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_14\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_6\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_14\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_12\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_13\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_6\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_0\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_1\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_6\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_6\ : std_logic;
signal \PWMInstance7.periodCounterZ0Z_7\ : std_logic;
signal \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_6\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_8\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_13\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_11\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_12\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_5\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_4\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_7\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_6\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_15\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_1\ : std_logic;
signal \PWMInstance7.PWMPulseWidthCountZ0Z_0\ : std_logic;
signal \PWMInstance7.pwmWrite_0_7\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_9\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_8\ : std_logic;
signal \RST_c_i\ : std_logic;
signal \ch0_B_c\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_2\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_3\ : std_logic;
signal \PWMInstance1.un1_periodCounter12_1_0_a2_0_0_cascade_\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_4\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_0\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_1\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_7\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_8\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_5\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_9\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_6\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_14\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_15\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_11\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_13\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_0\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_1\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_2\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_3\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_4\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_5\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_6\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_7\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_8\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_9\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_10\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_11\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_12\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_13\ : std_logic;
signal \QuadInstance2.un1_Quad_cry_14\ : std_logic;
signal \QuadInstance2.Quad_RNI8TLE2Z0Z_9\ : std_logic;
signal \QuadInstance2.Quad_RNIHU2G2Z0Z_11\ : std_logic;
signal \QuadInstance2.Quad_RNI0LLE2Z0Z_1\ : std_logic;
signal \QuadInstance2.Quad_RNIGT2G2Z0Z_10\ : std_logic;
signal \QuadInstance2.Quad_RNIIV2G2Z0Z_12\ : std_logic;
signal \QuadInstance2.Quad_RNI6RLE2Z0Z_7\ : std_logic;
signal \QuadInstance2.Quad_RNI7SLE2Z0Z_8\ : std_logic;
signal \QuadInstance2.Quad_RNI3OLE2Z0Z_4\ : std_logic;
signal \QuadInstance2.un1_Quad_axb_15\ : std_logic;
signal \QuadInstance2.count_enable_cascade_\ : std_logic;
signal \QuadInstance2.Quad_RNI1MLE2Z0Z_2\ : std_logic;
signal \QuadInstance2.un1_count_enable_i_a2_0_1_cascade_\ : std_logic;
signal \QuadInstance2.Quad_RNI2NLE2Z0Z_3\ : std_logic;
signal \QuadInstance2.Quad_RNI4PLE2Z0Z_5\ : std_logic;
signal \QuadInstance2.Quad_RNI5QLE2Z0Z_6\ : std_logic;
signal \QuadInstance2.delayedCh_AZ0Z_1\ : std_logic;
signal \QuadInstance2.delayedCh_AZ0Z_2\ : std_logic;
signal \QuadInstance2.Quad_RNIK13G2Z0Z_14\ : std_logic;
signal \QuadInstance2.delayedCh_BZ0Z_1\ : std_logic;
signal \QuadInstance2.delayedCh_BZ0Z_2\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_0\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_0\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_0\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_0\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_1\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_0\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_2\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_0\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_3\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_0\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_4\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_0\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_5\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_0\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_6\ : std_logic;
signal \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_7\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \PWM1_c\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_2\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_3\ : std_logic;
signal \PWMInstance0.un1_periodCounter12_1_0_a2_0_0_cascade_\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_5\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_4\ : std_logic;
signal \pwmWrite_fastZ0Z_0\ : std_logic;
signal \PWMInstance0.clkCountZ0Z_1\ : std_logic;
signal \PWMInstance0.clkCountZ0Z_0\ : std_logic;
signal \PWMInstance0.periodCounter12_cascade_\ : std_logic;
signal \PWMInstance0.un1_periodCounter12_1_0_a2_0_6\ : std_logic;
signal \PWMInstance0.un1_periodCounter12_1_0_a2_0_10\ : std_logic;
signal \PWMInstance0.un1_periodCounter12_1_0_a2_0_14_cascade_\ : std_logic;
signal \PWMInstance0.un1_periodCounter12_1_0_a2_0_12\ : std_logic;
signal \PWMInstance0.periodCounter12\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_0\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_2\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_1\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_3\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_2\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_4\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_3\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_5\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_4\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_5\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_6\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_7\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_8\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_9\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_10\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_11\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_12\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_13\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_14\ : std_logic;
signal \PWMInstance0.un1_periodCounter_2_cry_15\ : std_logic;
signal \bfn_7_18_0_\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_16\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_0\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_0\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_2\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_1\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_3\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_2\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_4\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_3\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_5\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_4\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_6\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_5\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_6\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_7\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_8\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_9\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_8\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_10\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_9\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_11\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_10\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_12\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_11\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_13\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_12\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_14\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_13\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_14\ : std_logic;
signal \PWMInstance1.un1_periodCounter_2_cry_15\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_0\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_1\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_2\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_4\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_3\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_4\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_5\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_6\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_7\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \PWM5_c\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_12\ : std_logic;
signal \PWMInstance1.PWMPulseWidthCountZ0Z_10\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_9\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_10\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_14\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_12\ : std_logic;
signal \QuadInstance7.un1_count_enable_i_a2_0_1_cascade_\ : std_logic;
signal \QuadInstance7.count_enable_cascade_\ : std_logic;
signal \QuadInstance7.un1_count_enable_i_a2_0_1\ : std_logic;
signal \QuadInstance7.delayedCh_AZ0Z_1\ : std_logic;
signal \QuadInstance7.delayedCh_AZ0Z_2\ : std_logic;
signal \QuadInstance7.delayedCh_BZ0Z_1\ : std_logic;
signal \QuadInstance7.delayedCh_BZ0Z_2\ : std_logic;
signal \PWMInstance1.un1_periodCounter12_1_0_a2_0\ : std_logic;
signal \PWMInstance1.pwmWrite_0_1\ : std_logic;
signal \pwmWriteZ0Z_1\ : std_logic;
signal \PWMInstance1.clkCountZ0Z_1\ : std_logic;
signal \PWMInstance1.clkCountZ0Z_0\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_16\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_7\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_15\ : std_logic;
signal \PWMInstance1.periodCounterZ0Z_1\ : std_logic;
signal \PWMInstance1.un1_periodCounter12_1_0_a2_0_6_cascade_\ : std_logic;
signal \PWMInstance1.periodCounter12\ : std_logic;
signal \PWMInstance1.un1_periodCounter12_1_0_a2_0_10\ : std_logic;
signal \PWMInstance1.un1_periodCounter12_1_0_a2_0_9\ : std_logic;
signal \PWMInstance1.un1_periodCounter12_1_0_a2_0_14_cascade_\ : std_logic;
signal \PWMInstance1.un1_periodCounter12_1_0_a2_0_12\ : std_logic;
signal \PWMInstance1.out_0_sqmuxa\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_4\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_2\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_3\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_14\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_4\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_15\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_9\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_9\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_8\ : std_logic;
signal \pwmWriteZ0Z_0\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_12\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_4\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_6\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_7\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_15\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_14\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_14\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_15\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_10\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_11\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_10\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_11\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_13\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_12\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_12\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNOZ0\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_0\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNOZ0\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_1\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNOZ0\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_2\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNOZ0\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_3\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNOZ0\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_4\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNOZ0\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_5\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNOZ0\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_6\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_7\ : std_logic;
signal \PWMInstance0.un1_periodCounter12_1_0_a2_0\ : std_logic;
signal \PWMInstance0.out_0_sqmuxa\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \PWM0_c\ : std_logic;
signal \ch7_B_c\ : std_logic;
signal \QuadInstance7.delayedCh_BZ0Z_0\ : std_logic;
signal \PWM0_obufLegalizeSB_DFFNet\ : std_logic;
signal \PWM1_obufLegalizeSB_DFFNet\ : std_logic;
signal \PWM6_obufLegalizeSB_DFFNet\ : std_logic;
signal \PWM7_obufLegalizeSB_DFFNet\ : std_logic;
signal \ch3_B_c\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_4\ : std_logic;
signal \ch5_A_c\ : std_logic;
signal \QuadInstance5.delayedCh_AZ0Z_0\ : std_logic;
signal \QuadInstance5.un1_count_enable_i_a2_0_1_cascade_\ : std_logic;
signal \QuadInstance2.un1_count_enable_i_a2_0_1\ : std_logic;
signal \QuadInstance2.Quad_RNIJ03G2Z0Z_13\ : std_logic;
signal \QuadInstance5.un1_count_enable_i_a2_0_1\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \QuadInstance7.Quad_RNI85VV2Z0Z_1\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_0\ : std_logic;
signal \QuadInstance7.Quad_RNI96VV2Z0Z_2\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_1\ : std_logic;
signal \QuadInstance7.Quad_RNIA7VV2Z0Z_3\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_2\ : std_logic;
signal \QuadInstance7.Quad_RNIB8VV2Z0Z_4\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_3\ : std_logic;
signal \QuadInstance7.Quad_RNIC9VV2Z0Z_5\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_4\ : std_logic;
signal \QuadInstance7.Quad_RNIDAVV2Z0Z_6\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_5\ : std_logic;
signal \QuadInstance7.Quad_RNIEBVV2Z0Z_7\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_6\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_7\ : std_logic;
signal \QuadInstance7.Quad_RNIFCVV2Z0Z_8\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \QuadInstance7.Quad_RNIGDVV2Z0Z_9\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_8\ : std_logic;
signal \QuadInstance7.Quad_RNIOIKU2Z0Z_10\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_9\ : std_logic;
signal \QuadInstance7.Quad_RNIPJKU2Z0Z_11\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_11\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_10\ : std_logic;
signal \QuadInstance7.Quad_RNIQKKU2Z0Z_12\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_12\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_11\ : std_logic;
signal \QuadInstance7.Quad_RNIRLKU2Z0Z_13\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_12\ : std_logic;
signal \QuadInstance7.Quad_RNISMKU2Z0Z_14\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_13\ : std_logic;
signal \QuadInstance7.un1_Quad_axb_15\ : std_logic;
signal \QuadInstance7.un1_Quad_cry_14\ : std_logic;
signal \pwmWrite_fastZ0Z_1\ : std_logic;
signal \pwmWriteZ0Z_7\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_4\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_0\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_1\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_4\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_6\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_7\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_0\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_0\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_1\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_2\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_3\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_4\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_6\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_5\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_6\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_7\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_8\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_8\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_9\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_10\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_11\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_13\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_12\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_13\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_14\ : std_logic;
signal \PWMInstance5.un1_periodCounter_2_cry_15\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_8\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_6\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_13\ : std_logic;
signal \PWMInstance0.un1_periodCounter12_1_0_a2_0_9\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_0\ : std_logic;
signal \PWMInstance0.periodCounterZ0Z_1\ : std_logic;
signal \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNOZ0\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_0\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_1\ : std_logic;
signal \PWMInstance0.PWMPulseWidthCountZ0Z_7\ : std_logic;
signal \PWMInstance0.pwmWrite_0_0\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_13\ : std_logic;
signal \ch5_B_c\ : std_logic;
signal \QuadInstance5.delayedCh_BZ0Z_0\ : std_logic;
signal \QuadInstance2.count_enable\ : std_logic;
signal \QuadInstance5.delayedCh_BZ0Z_1\ : std_logic;
signal \QuadInstance5.delayedCh_AZ0Z_1\ : std_logic;
signal \QuadInstance5.delayedCh_AZ0Z_2\ : std_logic;
signal \QuadInstance5.delayedCh_BZ0Z_2\ : std_logic;
signal \QuadInstance5.count_enable_cascade_\ : std_logic;
signal \QuadInstance5.count_enable\ : std_logic;
signal \bfn_10_6_0_\ : std_logic;
signal \QuadInstance5.Quad_RNIOUKI2Z0Z_1\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_4_1\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_0\ : std_logic;
signal \QuadInstance5.Quad_RNIPVKI2Z0Z_2\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_1\ : std_logic;
signal \QuadInstance5.Quad_RNIQ0LI2Z0Z_3\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_2\ : std_logic;
signal \QuadInstance5.Quad_RNIR1LI2Z0Z_4\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_3\ : std_logic;
signal \QuadInstance5.Quad_RNIS2LI2Z0Z_5\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_4\ : std_logic;
signal \QuadInstance5.Quad_RNIT3LI2Z0Z_6\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_5\ : std_logic;
signal \QuadInstance5.Quad_RNIU4LI2Z0Z_7\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_6\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_7\ : std_logic;
signal \QuadInstance5.Quad_RNIV5LI2Z0Z_8\ : std_logic;
signal \bfn_10_7_0_\ : std_logic;
signal \QuadInstance5.Quad_RNI07LI2Z0Z_9\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_8\ : std_logic;
signal \QuadInstance5.Quad_RNI8AQ82Z0Z_10\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_9\ : std_logic;
signal \QuadInstance5.Quad_RNI9BQ82Z0Z_11\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_10\ : std_logic;
signal \QuadInstance5.Quad_RNIACQ82Z0Z_12\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_12\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_11\ : std_logic;
signal \QuadInstance5.Quad_RNIBDQ82Z0Z_13\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_13\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_12\ : std_logic;
signal \QuadInstance5.Quad_RNICEQ82Z0Z_14\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_14\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_13\ : std_logic;
signal \QuadInstance5.un1_Quad_axb_15\ : std_logic;
signal \QuadInstance5.un1_Quad_cry_14\ : std_logic;
signal \bfn_10_8_0_\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_0\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_1\ : std_logic;
signal \QuadInstance3.Quad_RNIAQAL1Z0Z_3\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_2\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_3\ : std_logic;
signal \QuadInstance3.Quad_RNICSAL1Z0Z_5\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_4\ : std_logic;
signal \QuadInstance3.Quad_RNIDTAL1Z0Z_6\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_5\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_6\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_7\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_8\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_9\ : std_logic;
signal \QuadInstance3.Quad_RNIP20J1Z0Z_11\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_10\ : std_logic;
signal \QuadInstance3.Quad_RNIQ30J1Z0Z_12\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_11\ : std_logic;
signal \QuadInstance3.Quad_RNIR40J1Z0Z_13\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_12\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_13\ : std_logic;
signal \QuadInstance3.un1_Quad_cry_14\ : std_logic;
signal \QuadInstance3.count_enable_cascade_\ : std_logic;
signal \QuadInstance3.Quad_RNI8OAL1Z0Z_1\ : std_logic;
signal \QuadInstance3.un1_count_enable_i_a2_0_1_cascade_\ : std_logic;
signal \QuadInstance3.Quad_RNI9PAL1Z0Z_2\ : std_logic;
signal \QuadInstance3.Quad_RNIO10J1Z0Z_10\ : std_logic;
signal \QuadInstance3.Quad_RNIFVAL1Z0Z_8\ : std_logic;
signal \QuadInstance3.Quad_RNIG0BL1Z0Z_9\ : std_logic;
signal \QuadInstance3.Quad_RNIBRAL1Z0Z_4\ : std_logic;
signal \QuadInstance3.Quad_RNIS50J1Z0Z_14\ : std_logic;
signal \QuadInstance3.delayedCh_BZ0Z_2\ : std_logic;
signal \QuadInstance3.delayedCh_AZ0Z_2\ : std_logic;
signal \QuadInstance3.delayedCh_AZ0Z_1\ : std_logic;
signal \QuadInstance3.Quad_RNIEUAL1Z0Z_7\ : std_logic;
signal \QuadInstance3.un1_count_enable_i_a2_0_1\ : std_logic;
signal \QuadInstance3.count_enable\ : std_logic;
signal \QuadInstance3.un1_Quad_axb_15\ : std_logic;
signal \QuadInstance3.delayedCh_BZ0Z_0\ : std_logic;
signal \QuadInstance3.delayedCh_BZ0Z_1\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_4\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_2\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_14\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_12\ : std_logic;
signal \PWMInstance5.un1_periodCounter12_1_0_a2_0_0_cascade_\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_4\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_4\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_5\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_10\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_10\ : std_logic;
signal \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_4\ : std_logic;
signal \PWMInstance5.PWMPulseWidthCountZ0Z_11\ : std_logic;
signal \PWMInstance5.un1_periodCounter12_1_0_a2_0\ : std_logic;
signal \PWMInstance5.pwmWrite_0_5\ : std_logic;
signal \PWMInstance5.clkCountZ0Z_1\ : std_logic;
signal \PWMInstance5.clkCountZ0Z_0\ : std_logic;
signal \PWMInstance5.periodCounter12\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_15\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_1\ : std_logic;
signal \PWMInstance5.periodCounter12_cascade_\ : std_logic;
signal \PWMInstance5.un1_periodCounter12_1_0_a2_0_9\ : std_logic;
signal \PWMInstance5.un1_periodCounter12_1_0_a2_0_14_cascade_\ : std_logic;
signal \PWMInstance5.un1_periodCounter12_1_0_a2_0_12\ : std_logic;
signal \PWMInstance5.out_0_sqmuxa\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_9\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_5\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_11\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_3\ : std_logic;
signal \PWMInstance5.un1_periodCounter12_1_0_a2_0_10\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_16\ : std_logic;
signal \PWMInstance5.periodCounterZ0Z_7\ : std_logic;
signal \PWMInstance5.un1_periodCounter12_1_0_a2_0_6\ : std_logic;
signal \PWMInstance6.un1_periodCounter12_1_0_a2_0_0_cascade_\ : std_logic;
signal \PWMInstance6.un1_periodCounter12_1_0_a2_0_12_cascade_\ : std_logic;
signal \PWMInstance6.un1_periodCounter12_1_0_a2_0_10\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_2\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_3\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_4\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_2\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_2\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_6\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_2\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_3\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_4\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_6\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_6\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_9\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_8\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_3\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_7\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_7\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_7\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_5\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_7\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_11\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_10\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_11\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_8\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_9\ : std_logic;
signal \dataRead5_13\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_13\ : std_logic;
signal \dataRead2_13\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_13\ : std_logic;
signal \dataRead3_13\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_12\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_8\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_14\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_2\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_14\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_10\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_11\ : std_logic;
signal \OutReg_ess_RNO_2Z0Z_13\ : std_logic;
signal \dataRead5_11\ : std_logic;
signal \OutReg_0_5_i_m3_i_m3_ns_1_11_cascade_\ : std_logic;
signal \dataRead3_14\ : std_logic;
signal \dataRead2_14\ : std_logic;
signal \dataRead7_14\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_14_cascade_\ : std_logic;
signal \pwmWrite_fastZ0Z_5\ : std_logic;
signal \pwmWriteZ0Z_5\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_0\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_2\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_1\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_3\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_2\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_4\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_3\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_5\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_4\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_5\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_6\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_7\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_8\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_9\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_10\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_11\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_12\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_13\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_14\ : std_logic;
signal \PWMInstance6.un1_periodCounter_2_cry_15\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \ch3_A_c\ : std_logic;
signal \QuadInstance3.delayedCh_AZ0Z_0\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_2_5\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_5\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_5\ : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_0\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_2\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_1\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_3\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_2\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_3\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_5\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_4\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_6\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_5\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_7\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_6\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_7\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_8\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_8\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_9\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_11\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_10\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_12\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_11\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_13\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_12\ : std_logic;
signal \QuadInstance6.Quad_RNIKINB1Z0Z_14\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_13\ : std_logic;
signal \QuadInstance6.un1_Quad_axb_15\ : std_logic;
signal \QuadInstance6.un1_Quad_cry_14\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_5_1\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_8\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_14\ : std_logic;
signal \dataRead6_14\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_10\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_10\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_9\ : std_logic;
signal \QuadInstance6.Quad_RNI02A91Z0Z_1\ : std_logic;
signal \QuadInstance6.count_enable_cascade_\ : std_logic;
signal \QuadInstance6.Quad_RNI13A91Z0Z_2\ : std_logic;
signal \QuadInstance6.Quad_RNIHFNB1Z0Z_11\ : std_logic;
signal \QuadInstance6.Quad_RNI24A91Z0Z_3\ : std_logic;
signal \QuadInstance6.Quad_RNI46A91Z0Z_5\ : std_logic;
signal \QuadInstance6.Quad_RNI8AA91Z0Z_9\ : std_logic;
signal \QuadInstance6.Quad_RNI79A91Z0Z_8\ : std_logic;
signal \QuadInstance6.un1_count_enable_i_a2_0_1_cascade_\ : std_logic;
signal \QuadInstance6.Quad_RNI35A91Z0Z_4\ : std_logic;
signal \QuadInstance6.Quad_RNIIGNB1Z0Z_12\ : std_logic;
signal \QuadInstance6.Quad_RNI57A91Z0Z_6\ : std_logic;
signal \QuadInstance6.Quad_RNI68A91Z0Z_7\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_13\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_13\ : std_logic;
signal \dataRead7_11\ : std_logic;
signal \dataRead6_11\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_11_cascade_\ : std_logic;
signal \OutReg_ess_RNO_2Z0Z_11\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_11_cascade_\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_13\ : std_logic;
signal \data_receivedZ0Z_18\ : std_logic;
signal \data_receivedZ0Z_17\ : std_logic;
signal \data_receivedZ0Z_16\ : std_logic;
signal \data_receivedZ0Z_15\ : std_logic;
signal \PWMInstance6.clkCountZ0Z_0\ : std_logic;
signal \PWMInstance6.clkCountZ0Z_1\ : std_logic;
signal \pwmWrite_fastZ0Z_6\ : std_logic;
signal \pwmWriteZ0Z_6\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_16\ : std_logic;
signal \PWMInstance6.un1_periodCounter12_1_0_a2_0_6_cascade_\ : std_logic;
signal \PWMInstance6.periodCounter12\ : std_logic;
signal \PWMInstance6.un1_periodCounter12_1_0_a2_0_14\ : std_logic;
signal \ch6_A_c\ : std_logic;
signal \QuadInstance6.delayedCh_AZ0Z_0\ : std_logic;
signal \PWMInstance6.un1_periodCounter12_1_0_a2_0_9\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_0\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_1\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_0\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_1\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_6\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_7\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_6\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_7\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_8\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_9\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_5\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_5\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_0\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_5\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_1\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_5\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_2\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_5\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_3\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_4\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_5\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_6\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_7\ : std_logic;
signal \PWMInstance6.un1_periodCounter12_1_0_a2_0\ : std_logic;
signal \PWMInstance6.out_0_sqmuxa\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \PWM6_c\ : std_logic;
signal \PWM5_obufLegalizeSB_DFFNet\ : std_logic;
signal \ch2_A_c\ : std_logic;
signal \QuadInstance2.delayedCh_AZ0Z_0\ : std_logic;
signal \dataRead5_4\ : std_logic;
signal \OutReg_ess_RNO_2Z0Z_4_cascade_\ : std_logic;
signal \dataRead2_4\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_4_cascade_\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_4\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_4\ : std_logic;
signal \ch0_A_c\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_6\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_4\ : std_logic;
signal \dataRead6_4\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_4\ : std_logic;
signal \dataRead7_4\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_0_1\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_0\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_2\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_1\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_3\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_2\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_4\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_3\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_5\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_4\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_6\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_5\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_7\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_6\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_7\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_8\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_8\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_10\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_9\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_11\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_10\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_11\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_12\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_14\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_13\ : std_logic;
signal \QuadInstance1.un1_Quad_cry_14\ : std_logic;
signal \QuadInstance6.Quad_RNO_0_6_9\ : std_logic;
signal \QuadInstance2.Quad_RNO_0_1_1\ : std_logic;
signal \quadWriteZ0Z_2\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_2_1\ : std_logic;
signal \quadWriteZ0Z_3\ : std_logic;
signal \QuadInstance3.Quad_RNO_0_3_4\ : std_logic;
signal \dataRead3_4\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_9\ : std_logic;
signal \QuadInstance7.count_enable\ : std_logic;
signal \QuadInstance6.delayedCh_BZ0Z_2\ : std_logic;
signal \QuadInstance6.Quad_RNIGENB1Z0Z_10\ : std_logic;
signal \QuadInstance6.delayedCh_AZ0Z_1\ : std_logic;
signal \QuadInstance6.delayedCh_AZ0Z_2\ : std_logic;
signal \dataRead6_13\ : std_logic;
signal \quadWriteZ0Z_6\ : std_logic;
signal \QuadInstance6.un1_count_enable_i_a2_0_1\ : std_logic;
signal \QuadInstance6.count_enable\ : std_logic;
signal \QuadInstance6.Quad_RNIJHNB1Z0Z_13\ : std_logic;
signal \QuadInstance6.delayedCh_BZ0Z_1\ : std_logic;
signal \dataRead2_11\ : std_logic;
signal \dataRead3_11\ : std_logic;
signal \OutReg_0_4_i_m3_i_m3_ns_1_11\ : std_logic;
signal \dataRead5_12\ : std_logic;
signal \dataRead2_12\ : std_logic;
signal \dataRead3_12\ : std_logic;
signal \dataRead6_12\ : std_logic;
signal \dataRead7_12\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_12_cascade_\ : std_logic;
signal \OutReg_esr_RNO_1Z0Z_12_cascade_\ : std_logic;
signal \OutReg_esr_RNO_2Z0Z_12\ : std_logic;
signal \OutRegZ0Z_11\ : std_logic;
signal \OutReg_esr_RNO_0Z0Z_12_cascade_\ : std_logic;
signal \OutRegZ0Z_12\ : std_logic;
signal \data_receivedZ0Z_12\ : std_logic;
signal \data_receivedZ0Z_13\ : std_logic;
signal \data_receivedZ0Z_14\ : std_logic;
signal \data_receivedZ0Z_10\ : std_logic;
signal \data_receivedZ0Z_11\ : std_logic;
signal \data_received_esr_RNIMIH31Z0Z_19_cascade_\ : std_logic;
signal \data_receivedZ0Z_19\ : std_logic;
signal \data_receivedZ0Z_23\ : std_logic;
signal \data_received_esr_RNIMIH31_0Z0Z_19_cascade_\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_5\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_8\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_15\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_14\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_5\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_14\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_15\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_10\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_11\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_11\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_5\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_10\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_13\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_12\ : std_logic;
signal \PWMInstance6.periodCounterZ0Z_13\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_12\ : std_logic;
signal \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_5\ : std_logic;
signal \PWMInstance4.un1_periodCounter12_1_0_a2_0_0_cascade_\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_4\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_5\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_10\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_11\ : std_logic;
signal \ch2_B_c\ : std_logic;
signal \QuadInstance2.delayedCh_BZ0Z_0\ : std_logic;
signal \ch4_B_c\ : std_logic;
signal \ch4_A_c\ : std_logic;
signal \dataRead1_4\ : std_logic;
signal \QuadInstance1.Quad_RNIRK0OZ0Z_4\ : std_logic;
signal \QuadInstance1.delayedCh_BZ0Z_1\ : std_logic;
signal \QuadInstance1.count_enable_cascade_\ : std_logic;
signal \QuadInstance1.Quad_RNIOH0OZ0Z_1\ : std_logic;
signal \QuadInstance1.Quad_RNITM0OZ0Z_6\ : std_logic;
signal \QuadInstance1.Quad_RNISL0OZ0Z_5\ : std_logic;
signal \QuadInstance1.delayedCh_AZ0Z_2\ : std_logic;
signal \QuadInstance1.delayedCh_BZ0Z_2\ : std_logic;
signal \QuadInstance1.delayedCh_AZ0Z_1\ : std_logic;
signal \QuadInstance1.Quad_RNI0Q0OZ0Z_9\ : std_logic;
signal \QuadInstance1.Quad_RNI8P5DZ0Z_10\ : std_logic;
signal \data_received_esr_RNIMIH31Z0Z_19\ : std_logic;
signal \dataRead1_11\ : std_logic;
signal \QuadInstance1.Quad_RNI9Q5DZ0Z_11\ : std_logic;
signal \dataRead3_5\ : std_logic;
signal \dataRead2_5\ : std_logic;
signal \QuadInstance1.Quad_RNIUN0OZ0Z_7\ : std_logic;
signal \QuadInstance1.Quad_RNIPI0OZ0Z_2\ : std_logic;
signal \QuadInstance1.Quad_RNIQJ0OZ0Z_3\ : std_logic;
signal \QuadInstance1.Quad_RNIAR5DZ0Z_12\ : std_logic;
signal \QuadInstance1.Quad_RNIBS5DZ0Z_13\ : std_logic;
signal \QuadInstance1.Quad_RNICT5DZ0Z_14\ : std_logic;
signal \QuadInstance1.Quad_RNIVO0OZ0Z_8\ : std_logic;
signal \QuadInstance1.un1_count_enable_i_a2_0_1\ : std_logic;
signal \QuadInstance1.un1_Quad_axb_15\ : std_logic;
signal \QuadInstance1.count_enable\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_12\ : std_logic;
signal \dataRead1_12\ : std_logic;
signal \quadWriteZ0Z_1\ : std_logic;
signal \QuadInstance1.Quad_RNO_0_1_13\ : std_logic;
signal \dataRead1_13\ : std_logic;
signal \dataRead1_1\ : std_logic;
signal \dataRead5_1\ : std_logic;
signal \OutReg_ess_RNO_2Z0Z_1_cascade_\ : std_logic;
signal \dataRead2_1\ : std_logic;
signal \dataRead3_1\ : std_logic;
signal \dataRead6_1\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_1_cascade_\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_1\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_1\ : std_logic;
signal \dataRead2_3\ : std_logic;
signal \dataRead3_3\ : std_logic;
signal \dataRead3_15\ : std_logic;
signal \dataRead2_15\ : std_logic;
signal \dataRead7_15\ : std_logic;
signal \dataRead6_15\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_15_cascade_\ : std_logic;
signal \dataRead5_15\ : std_logic;
signal \dataRead1_15\ : std_logic;
signal \data_receivedZ0Z_5\ : std_logic;
signal \data_receivedZ0Z_6\ : std_logic;
signal \data_receivedZ0Z_7\ : std_logic;
signal \data_receivedZ0Z_8\ : std_logic;
signal \data_receivedZ0Z_9\ : std_logic;
signal \N_870_i\ : std_logic;
signal \pwmWriteZ0Z_3\ : std_logic;
signal \pwmWrite_fastZ0Z_3\ : std_logic;
signal \PWMInstance3.clkCountZ0Z_1\ : std_logic;
signal \PWMInstance3.clkCountZ0Z_0\ : std_logic;
signal \PWMInstance3.un1_periodCounter12_1_0_a2_0_6_cascade_\ : std_logic;
signal \PWMInstance3.un1_periodCounter12_1_0_a2_0_14_cascade_\ : std_logic;
signal \PWMInstance6.PWMPulseWidthCountZ0Z_9\ : std_logic;
signal \PWMInstance6.pwmWrite_0_6\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_3\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_2\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_14\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_15\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_12\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_13\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_0\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_2\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_1\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_3\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_2\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_4\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_3\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_5\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_4\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_5\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_6\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_7\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_8\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_10\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_9\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_11\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_10\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_12\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_11\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_12\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_14\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_13\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_14\ : std_logic;
signal \PWMInstance4.un1_periodCounter_2_cry_15\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \bfn_15_1_0_\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_3\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_0\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_3\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_1\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_2\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_3\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_3\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_4\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_3\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_5\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_3\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_6\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_7\ : std_logic;
signal \bfn_15_2_0_\ : std_logic;
signal \PWM4_c\ : std_logic;
signal \bfn_15_3_0_\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_3_1\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_0\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_1\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_2\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_4\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_3\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_4\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_5\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_6\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_7\ : std_logic;
signal \bfn_15_4_0_\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_9\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_8\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_9\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_10\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_11\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_12\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_13\ : std_logic;
signal \QuadInstance4.un1_Quad_axb_15\ : std_logic;
signal \QuadInstance4.un1_Quad_cry_14\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_6\ : std_logic;
signal \QuadInstance4.Quad_RNIL00S1Z0Z_6\ : std_logic;
signal \QuadInstance4.Quad_RNI06TL1Z0Z_10\ : std_logic;
signal \QuadInstance4.Quad_RNI17TL1Z0Z_11\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_11\ : std_logic;
signal \dataRead4_11\ : std_logic;
signal \dataRead4_6\ : std_logic;
signal \dataRead1_6\ : std_logic;
signal \dataRead5_6\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_6_cascade_\ : std_logic;
signal \QuadInstance4.Quad_RNIO30S1Z0Z_9\ : std_logic;
signal \QuadInstance4.Quad_RNIM10S1Z0Z_7\ : std_logic;
signal \dataRead4_15\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_15\ : std_logic;
signal \dataRead1_9\ : std_logic;
signal \dataRead5_9\ : std_logic;
signal \OutReg_ess_RNO_2Z0Z_9_cascade_\ : std_logic;
signal \dataRead3_9\ : std_logic;
signal \dataRead2_9\ : std_logic;
signal \dataRead6_9\ : std_logic;
signal \dataRead7_9\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_9_cascade_\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_9\ : std_logic;
signal \dataRead4_9\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_9\ : std_logic;
signal \N_45_0_g\ : std_logic;
signal \N_1187_g\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_13\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_13\ : std_logic;
signal \dataRead7_13\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_3\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_7_3\ : std_logic;
signal \quadWriteZ0Z_7\ : std_logic;
signal \QuadInstance7.Quad_RNO_0_6_1\ : std_logic;
signal \dataRead7_1\ : std_logic;
signal \quadWriteZ0Z_5\ : std_logic;
signal \QuadInstance5.Quad_RNO_0_5_3\ : std_logic;
signal \GB_BUFFER_RST_c_i_g_THRU_CO\ : std_logic;
signal \dataRead5_7\ : std_logic;
signal \dataRead1_7\ : std_logic;
signal \OutReg_ess_RNO_2Z0Z_7_cascade_\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_7_cascade_\ : std_logic;
signal \dataRead2_7\ : std_logic;
signal \dataRead3_7\ : std_logic;
signal \dataRead6_7\ : std_logic;
signal \dataRead7_7\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_7_cascade_\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_7\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_9\ : std_logic;
signal \OutRegZ0Z_13\ : std_logic;
signal \OutRegZ0Z_14\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_5\ : std_logic;
signal \PWMInstance3.un1_periodCounter12_1_0_a2_0_0_cascade_\ : std_logic;
signal \PWMInstance3.un1_periodCounter12_1_0_a2_0_12\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_4\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_11\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_10\ : std_logic;
signal \PWMInstance3.periodCounter12\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_0\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_1\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_2\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_4\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_3\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_4\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_5\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_6\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_7\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_8\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_10\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_9\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_10\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_11\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_12\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_13\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_14\ : std_logic;
signal \PWMInstance3.un1_periodCounter_2_cry_15\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_16\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_13\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_0\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_0\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_3\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_1\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_6\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_3\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_6\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_7\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_9\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_8\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_9\ : std_logic;
signal \PWMInstance4.PWMPulseWidthCountZ0Z_8\ : std_logic;
signal \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_3\ : std_logic;
signal \PWMInstance4.un1_periodCounter12_1_0_a2_0\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_16\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_7\ : std_logic;
signal \pwmWriteZ0Z_4\ : std_logic;
signal \PWMInstance4.pwmWrite_0_4\ : std_logic;
signal \pwmWrite_fastZ0Z_4\ : std_logic;
signal \PWMInstance4.clkCountZ0Z_1\ : std_logic;
signal \PWMInstance4.clkCountZ0Z_0\ : std_logic;
signal \PWMInstance4.periodCounter12\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_15\ : std_logic;
signal \PWMInstance4.periodCounterZ0Z_1\ : std_logic;
signal \PWMInstance4.periodCounter12_cascade_\ : std_logic;
signal \PWMInstance4.un1_periodCounter12_1_0_a2_0_6\ : std_logic;
signal \PWMInstance4.un1_periodCounter12_1_0_a2_0_10\ : std_logic;
signal \PWMInstance4.un1_periodCounter12_1_0_a2_0_9\ : std_logic;
signal \PWMInstance4.un1_periodCounter12_1_0_a2_0_14_cascade_\ : std_logic;
signal \PWMInstance4.un1_periodCounter12_1_0_a2_0_12\ : std_logic;
signal \PWMInstance4.out_0_sqmuxa\ : std_logic;
signal \ch6_B_c\ : std_logic;
signal \QuadInstance6.delayedCh_BZ0Z_0\ : std_logic;
signal \PWM4_obufLegalizeSB_DFFNet\ : std_logic;
signal \ch1_B_c\ : std_logic;
signal \QuadInstance1.delayedCh_BZ0Z_0\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_5\ : std_logic;
signal \dataRead4_5\ : std_logic;
signal \QuadInstance4.Quad_RNIKVVR1Z0Z_5\ : std_logic;
signal \QuadInstance4.Quad_RNI28TL1Z0Z_12\ : std_logic;
signal \QuadInstance4.count_enable_cascade_\ : std_logic;
signal \QuadInstance4.Quad_RNIHSVR1Z0Z_2\ : std_logic;
signal \dataRead4_1\ : std_logic;
signal \QuadInstance4.Quad_RNIGRVR1Z0Z_1\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_2\ : std_logic;
signal \dataRead4_2\ : std_logic;
signal \QuadInstance4.Quad_RNIITVR1Z0Z_3\ : std_logic;
signal \QuadInstance4.Quad_RNI39TL1Z0Z_13\ : std_logic;
signal \QuadInstance4.Quad_RNI4ATL1Z0Z_14\ : std_logic;
signal \QuadInstance4.delayedCh_BZ0Z_2\ : std_logic;
signal \dataRead4_4\ : std_logic;
signal \QuadInstance4.un1_count_enable_i_a2_0_1_cascade_\ : std_logic;
signal \QuadInstance4.Quad_RNIJUVR1Z0Z_4\ : std_logic;
signal \QuadInstance4.delayedCh_AZ0Z_0\ : std_logic;
signal \QuadInstance4.delayedCh_AZ0Z_1\ : std_logic;
signal \QuadInstance4.delayedCh_AZ0Z_2\ : std_logic;
signal \QuadInstance4.count_enable\ : std_logic;
signal \QuadInstance4.un1_count_enable_i_a2_0_1\ : std_logic;
signal \QuadInstance4.Quad_RNIN20S1Z0Z_8\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_8\ : std_logic;
signal \dataRead4_8\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_7\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_7\ : std_logic;
signal \dataRead4_7\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_12\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_12\ : std_logic;
signal \dataRead4_12\ : std_logic;
signal \dataRead4_13\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_13\ : std_logic;
signal \data_received_2_repZ0Z1\ : std_logic;
signal \dataRead4_3\ : std_logic;
signal \data_received_0_repZ0Z1\ : std_logic;
signal \dataRead5_3\ : std_logic;
signal \dataRead1_3\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_3_cascade_\ : std_logic;
signal \dataRead7_3\ : std_logic;
signal \dataRead6_3\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_3\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \OutReg_ess_RNO_2Z0Z_3\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \OutRegZ0Z_3\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_4\ : std_logic;
signal \dataRead6_6\ : std_logic;
signal \dataRead7_6\ : std_logic;
signal \OutReg_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \OutReg_esr_RNO_2Z0Z_6\ : std_logic;
signal \OutReg_esr_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \OutRegZ0Z_6\ : std_logic;
signal \dataRead2_6\ : std_logic;
signal \dataRead3_6\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_6\ : std_logic;
signal \dataRead5_14\ : std_logic;
signal \dataRead1_14\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_14_cascade_\ : std_logic;
signal \OutReg_esr_RNO_2Z0Z_14_cascade_\ : std_logic;
signal \OutReg_esr_RNO_1Z0Z_14\ : std_logic;
signal \OutReg_esr_RNO_0Z0Z_14\ : std_logic;
signal \dataWriteZ0Z_8\ : std_logic;
signal \dataWriteZ0Z_12\ : std_logic;
signal \dataWriteZ0Z_13\ : std_logic;
signal \dataWriteZ0Z_9\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_5\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_11\ : std_logic;
signal \PWMInstance3.un1_periodCounter12_1_0_a2_0_10\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_3\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_3\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_2\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_2\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_15\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_14\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_14\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_15\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_13\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_12\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_12\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_13\ : std_logic;
signal \PWMInstance3.un1_periodCounter12_1_0_a2_0_9\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_0\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_1\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_0\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_1\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_7\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_6\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_6\ : std_logic;
signal \dataWriteZ0Z_7\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_7\ : std_logic;
signal \PWMInstance3.pwmWrite_0_3\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_8\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_8\ : std_logic;
signal \PWMInstance3.periodCounterZ0Z_9\ : std_logic;
signal \PWMInstance3.PWMPulseWidthCountZ0Z_9\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_2\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_2\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_0\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_2\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_1\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_2\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_2\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_2\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_3\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_2\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_4\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_2\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_5\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_2\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_6\ : std_logic;
signal \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_7\ : std_logic;
signal \PWMInstance3.un1_periodCounter12_1_0_a2_0\ : std_logic;
signal \PWMInstance3.out_0_sqmuxa\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \PWM3_c\ : std_logic;
signal \ch7_A_c\ : std_logic;
signal \QuadInstance7.delayedCh_AZ0Z_0\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_10\ : std_logic;
signal \quadWriteZ0Z_4\ : std_logic;
signal \QuadInstance4.Quad_RNO_0_4_14\ : std_logic;
signal \dataRead4_14\ : std_logic;
signal \QuadInstance0.delayedCh_BZ0Z_0\ : std_logic;
signal \QuadInstance4.delayedCh_BZ0Z_0\ : std_logic;
signal \QuadInstance4.delayedCh_BZ0Z_1\ : std_logic;
signal \bfn_17_6_0_\ : std_logic;
signal \QuadInstance0.Quad_RNO_0Z0Z_1\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_0\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_2\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_1\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_3\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_2\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_4\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_3\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_5\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_4\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_6\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_5\ : std_logic;
signal \dataRead0_7\ : std_logic;
signal \QuadInstance0.Quad_RNIMKBH1Z0Z_7\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_7\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_6\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_7\ : std_logic;
signal \dataRead0_8\ : std_logic;
signal \QuadInstance0.Quad_RNINLBH1Z0Z_8\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_8\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \dataRead0_9\ : std_logic;
signal \QuadInstance0.Quad_RNIOMBH1Z0Z_9\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_9\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_8\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_9\ : std_logic;
signal \dataRead0_11\ : std_logic;
signal \QuadInstance0.Quad_RNI1M8Q1Z0Z_11\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_11\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_10\ : std_logic;
signal \dataRead0_12\ : std_logic;
signal \QuadInstance0.Quad_RNI2N8Q1Z0Z_12\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_12\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_11\ : std_logic;
signal \dataRead0_13\ : std_logic;
signal \QuadInstance0.Quad_RNI3O8Q1Z0Z_13\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_13\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_12\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_13\ : std_logic;
signal \QuadInstance0.un1_Quad_axb_15\ : std_logic;
signal \QuadInstance0.un1_Quad_cry_14\ : std_logic;
signal \dataRead0_15\ : std_logic;
signal \dataRead1_2\ : std_logic;
signal \dataRead5_2\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_2\ : std_logic;
signal \OutReg_esr_RNO_2Z0Z_2_cascade_\ : std_logic;
signal \OutReg_esr_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \OutRegZ0Z_2\ : std_logic;
signal \dataRead2_2\ : std_logic;
signal \dataRead3_2\ : std_logic;
signal \dataRead7_2\ : std_logic;
signal \dataRead6_2\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_2_cascade_\ : std_logic;
signal \OutReg_esr_RNO_1Z0Z_2\ : std_logic;
signal \dataRead0_0\ : std_logic;
signal \dataRead4_0\ : std_logic;
signal \dataRead1_0\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_0_cascade_\ : std_logic;
signal \dataRead5_0\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \dataRead3_0\ : std_logic;
signal \dataRead2_0\ : std_logic;
signal \dataRead6_0\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_0_cascade_\ : std_logic;
signal \dataRead7_0\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_0\ : std_logic;
signal \OutRegZ0Z_0\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_1\ : std_logic;
signal \OutRegZ0Z_1\ : std_logic;
signal \dataRead2_8\ : std_logic;
signal \dataRead3_8\ : std_logic;
signal \data_receivedZ0Z_3\ : std_logic;
signal \data_received_esr_RNI7L871Z0Z_3_cascade_\ : std_logic;
signal \OutReg_0_sqmuxa_0_a2_3_a2_2\ : std_logic;
signal \dataWriteZ0Z_0\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_0\ : std_logic;
signal \dataWriteZ0Z_1\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_1\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_7\ : std_logic;
signal \dataWriteZ0Z_6\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_6\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_8\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_9\ : std_logic;
signal \pwmWriteZ0Z_2\ : std_logic;
signal \pwmWrite_fastZ0Z_2\ : std_logic;
signal \PWMInstance2.clkCountZ0Z_1\ : std_logic;
signal \PWMInstance2.clkCountZ0Z_0\ : std_logic;
signal \PWMInstance2.un1_periodCounter12_1_0_a2_0_6_cascade_\ : std_logic;
signal \PWMInstance2.un1_periodCounter12_1_0_a2_0_9\ : std_logic;
signal \PWMInstance2.un1_periodCounter12_1_0_a2_0_14_cascade_\ : std_logic;
signal \PWMInstance2.un1_periodCounter12_1_0_a2_0_10\ : std_logic;
signal \dataWriteZ0Z_2\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_2\ : std_logic;
signal \dataWriteZ0Z_3\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_3\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_14\ : std_logic;
signal \dataWriteZ0Z_15\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_15\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_13\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_12\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_1\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_1\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_0\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_1\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_1\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_2\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_1\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_3\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_4\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_1\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_5\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_1\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_6\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_7\ : std_logic;
signal \PWMInstance2.un1_periodCounter12_1_0_a2_0\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \PWM2_c\ : std_logic;
signal \MOSI_c\ : std_logic;
signal \ch1_A_c\ : std_logic;
signal \QuadInstance1.delayedCh_AZ0Z_0\ : std_logic;
signal \QuadInstance0.delayedCh_AZ0Z_0\ : std_logic;
signal \data_received_0_repZ0Z2\ : std_logic;
signal \dataRead4_10\ : std_logic;
signal \data_received_2_repZ0Z2\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_10\ : std_logic;
signal \QuadInstance0.delayedCh_BZ0Z_1\ : std_logic;
signal \QuadInstance0.delayedCh_AZ0Z_2\ : std_logic;
signal \dataRead0_1\ : std_logic;
signal \QuadInstance0.count_enable_cascade_\ : std_logic;
signal \QuadInstance0.Quad_RNIGEBH1Z0Z_1\ : std_logic;
signal \dataRead0_10\ : std_logic;
signal \QuadInstance0.Quad_RNI0L8Q1Z0Z_10\ : std_logic;
signal \dataRead0_2\ : std_logic;
signal \QuadInstance0.Quad_RNIHFBH1Z0Z_2\ : std_logic;
signal \QuadInstance0.delayedCh_BZ0Z_2\ : std_logic;
signal \QuadInstance0.delayedCh_AZ0Z_1\ : std_logic;
signal \RST_c\ : std_logic;
signal \dataWriteZ0Z_14\ : std_logic;
signal \QuadInstance0.Quad_RNO_0_0_14\ : std_logic;
signal \dataRead0_14\ : std_logic;
signal \QuadInstance0.Quad_RNI4P8Q1Z0Z_14\ : std_logic;
signal \dataRead0_3\ : std_logic;
signal \QuadInstance0.Quad_RNIIGBH1Z0Z_3\ : std_logic;
signal \dataRead0_4\ : std_logic;
signal \QuadInstance0.Quad_RNIJHBH1Z0Z_4\ : std_logic;
signal \dataRead0_5\ : std_logic;
signal \QuadInstance0.Quad_RNIKIBH1Z0Z_5\ : std_logic;
signal \QuadInstance0.count_enable\ : std_logic;
signal \dataRead0_6\ : std_logic;
signal \QuadInstance0.un1_count_enable_i_a2_0_1\ : std_logic;
signal \QuadInstance0.Quad_RNILJBH1Z0Z_6\ : std_logic;
signal \data_receivedZ0Z_21\ : std_logic;
signal \data_receivedZ0Z_20\ : std_logic;
signal \data_receivedZ0Z_22\ : std_logic;
signal \data_received_esr_RNIMIH31_0Z0Z_19\ : std_logic;
signal \quadWriteZ0Z_0\ : std_logic;
signal \MOSIrZ0Z_0\ : std_logic;
signal \MOSIrZ0Z_1\ : std_logic;
signal \dataRead1_10\ : std_logic;
signal \dataRead5_10\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_10\ : std_logic;
signal \data_receivedZ0Z_4\ : std_logic;
signal \un1_OutReg51_4_0_i_o3_2_cascade_\ : std_logic;
signal \OutReg_21_m_0_a2_1_0\ : std_logic;
signal \OutReg_esr_RNO_2Z0Z_10\ : std_logic;
signal \OutRegZ0Z_9\ : std_logic;
signal \OutReg_esr_RNO_0Z0Z_10\ : std_logic;
signal \OutRegZ0Z_10\ : std_logic;
signal \data_received_fastZ0Z_2\ : std_logic;
signal \dataRead3_10\ : std_logic;
signal \data_received_fastZ0Z_0\ : std_logic;
signal \dataRead2_10\ : std_logic;
signal \dataRead7_10\ : std_logic;
signal \dataRead6_10\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_10_cascade_\ : std_logic;
signal \OutReg_esr_RNO_1Z0Z_10\ : std_logic;
signal \PWMInstance2.periodCounter12\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_0\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_1\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_0\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_1\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_3\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_2\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_3\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_4\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_6\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_5\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_7\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_6\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_7\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_8\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_9\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_8\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_9\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_10\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_11\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_13\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_12\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_13\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_15\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_14\ : std_logic;
signal \PWMInstance2.un1_periodCounter_2_cry_15\ : std_logic;
signal \PWMInstance2.out_0_sqmuxa\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_16\ : std_logic;
signal \PWMInstance0_N_42_g\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_5\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_1\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_14\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_2\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_4\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_12\ : std_logic;
signal \PWMInstance2.un1_periodCounter12_1_0_a2_0_0_cascade_\ : std_logic;
signal \PWMInstance2.un1_periodCounter12_1_0_a2_0_12\ : std_logic;
signal \dataWriteZ0Z_4\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_4\ : std_logic;
signal \dataWriteZ0Z_5\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_5\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_10\ : std_logic;
signal \PWMInstance2.periodCounterZ0Z_11\ : std_logic;
signal \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_1\ : std_logic;
signal \dataWriteZ0Z_10\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_10\ : std_logic;
signal \dataWriteZ0Z_11\ : std_logic;
signal \PWMInstance2.PWMPulseWidthCountZ0Z_11\ : std_logic;
signal \PWMInstance2.pwmWrite_0_2\ : std_logic;
signal \RST_c_i_g\ : std_logic;
signal \PWM2_obufLegalizeSB_DFFNet\ : std_logic;
signal \PWM3_obufLegalizeSB_DFFNet\ : std_logic;
signal \MISO_obufLegalizeSB_DFFNet\ : std_logic;
signal \internalOscilatorOutputNet\ : std_logic;
signal \dataRead5_5\ : std_logic;
signal \dataRead1_5\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_5\ : std_logic;
signal \dataRead6_5\ : std_logic;
signal \dataRead7_5\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_5\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_5_cascade_\ : std_logic;
signal \OutReg_ess_RNO_2Z0Z_5\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_5\ : std_logic;
signal \OutRegZ0Z_4\ : std_logic;
signal \OutRegZ0Z_5\ : std_logic;
signal \OutRegZ0Z_15\ : std_logic;
signal \dataOut_RNOZ0Z_0_cascade_\ : std_logic;
signal \MISO_c\ : std_logic;
signal \SSEL_c\ : std_logic;
signal \un1_bit_count_1_c1_cascade_\ : std_logic;
signal \OutReg_ess_RNO_1Z0Z_15\ : std_logic;
signal \OutReg_ess_RNO_2Z0Z_15\ : std_logic;
signal \OutReg_ess_RNO_0Z0Z_15\ : std_logic;
signal \bit_countZ0Z_0\ : std_logic;
signal \dataRead6_8\ : std_logic;
signal \data_receivedZ0Z_2\ : std_logic;
signal \dataRead7_8\ : std_logic;
signal \OutReg_0_4_i_m3_ns_1_8\ : std_logic;
signal \data_receivedZ0Z_1\ : std_logic;
signal \OutReg_esr_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \OutRegZ0Z_7\ : std_logic;
signal \OutReg_esr_RNO_0Z0Z_8_cascade_\ : std_logic;
signal \un1_OutReg51_4_0_i_o3_2\ : std_logic;
signal \OutRegZ0Z_8\ : std_logic;
signal \N_863_0\ : std_logic;
signal \OutReg_0_sqmuxa\ : std_logic;
signal \dataRead1_8\ : std_logic;
signal \dataRead5_8\ : std_logic;
signal \data_receivedZ0Z_0\ : std_logic;
signal \OutReg_0_5_i_m3_ns_1_8\ : std_logic;
signal \OutReg_esr_RNO_2Z0Z_8\ : std_logic;
signal \SSELrZ0Z_0\ : std_logic;
signal \SSELrZ0Z_2\ : std_logic;
signal \SCK_c\ : std_logic;
signal \bit_countZ0Z_2\ : std_logic;
signal \SCKr_RNIBA7CZ0Z_2\ : std_logic;
signal \SCKr_RNIBA7CZ0Z_2_cascade_\ : std_logic;
signal \N_45_0\ : std_logic;
signal \SCKrZ0Z_0\ : std_logic;
signal un1_bit_count_1_c1 : std_logic;
signal \bit_countZ0Z_1\ : std_logic;
signal \bit_count_RNIU615_0Z0Z_4\ : std_logic;
signal \bit_count_RNIU615_0Z0Z_4_cascade_\ : std_logic;
signal \SSELr_RNIGO0FZ0Z_1\ : std_logic;
signal \SSELrZ0Z_1\ : std_logic;
signal un1_bit_count_1_c3 : std_logic;
signal \bit_countZ0Z_3\ : std_logic;
signal \bit_countZ0Z_4\ : std_logic;
signal \un1_OutReg51_4_0_i_o3_3\ : std_logic;
signal \SCKrZ0Z_1\ : std_logic;
signal \SCKrZ0Z_2\ : std_logic;
signal myclk : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \PWM5_wire\ : std_logic;
signal \ch6_A_wire\ : std_logic;
signal \ch6_B_wire\ : std_logic;
signal \ch5_B_wire\ : std_logic;
signal \ch0_B_wire\ : std_logic;
signal \PWM6_wire\ : std_logic;
signal \PWM4_wire\ : std_logic;
signal \RST_wire\ : std_logic;
signal \MISO_wire\ : std_logic;
signal \ch5_A_wire\ : std_logic;
signal \ch2_B_wire\ : std_logic;
signal \ch4_B_wire\ : std_logic;
signal \PWM3_wire\ : std_logic;
signal \PWM1_wire\ : std_logic;
signal \ch4_A_wire\ : std_logic;
signal \ch7_A_wire\ : std_logic;
signal \ch3_B_wire\ : std_logic;
signal \PWM7_wire\ : std_logic;
signal \SCK_wire\ : std_logic;
signal \ch3_A_wire\ : std_logic;
signal \ch1_B_wire\ : std_logic;
signal \PWM2_wire\ : std_logic;
signal \MOSI_wire\ : std_logic;
signal \ch7_B_wire\ : std_logic;
signal \ch0_A_wire\ : std_logic;
signal \PWM0_wire\ : std_logic;
signal \SSEL_wire\ : std_logic;
signal \ch1_A_wire\ : std_logic;
signal \ch2_A_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    PWM5 <= \PWM5_wire\;
    \ch6_A_wire\ <= ch6_A;
    \ch6_B_wire\ <= ch6_B;
    \ch5_B_wire\ <= ch5_B;
    \ch0_B_wire\ <= ch0_B;
    PWM6 <= \PWM6_wire\;
    PWM4 <= \PWM4_wire\;
    \RST_wire\ <= RST;
    MISO <= \MISO_wire\;
    \ch5_A_wire\ <= ch5_A;
    \ch2_B_wire\ <= ch2_B;
    \ch4_B_wire\ <= ch4_B;
    PWM3 <= \PWM3_wire\;
    PWM1 <= \PWM1_wire\;
    \ch4_A_wire\ <= ch4_A;
    \ch7_A_wire\ <= ch7_A;
    \ch3_B_wire\ <= ch3_B;
    PWM7 <= \PWM7_wire\;
    \SCK_wire\ <= SCK;
    \ch3_A_wire\ <= ch3_A;
    \ch1_B_wire\ <= ch1_B;
    PWM2 <= \PWM2_wire\;
    \MOSI_wire\ <= MOSI;
    \ch7_B_wire\ <= ch7_B;
    \ch0_A_wire\ <= ch0_A;
    PWM0 <= \PWM0_wire\;
    \SSEL_wire\ <= SSEL;
    \ch1_A_wire\ <= ch1_A;
    \ch2_A_wire\ <= ch2_A;

    \CLK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39370\,
            DIN => \N__39369\,
            DOUT => \N__39368\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39370\,
            PADOUT => \N__39369\,
            PADIN => \N__39368\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWM5_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39361\,
            DIN => \N__39360\,
            DOUT => \N__39359\,
            PACKAGEPIN => \PWM5_wire\
        );

    \PWM5_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39361\,
            PADOUT => \N__39360\,
            PADIN => \N__39359\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__21357\,
            DIN0 => OPEN,
            DOUT0 => \N__16401\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch6_A_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39352\,
            DIN => \N__39351\,
            DOUT => \N__39350\,
            PACKAGEPIN => \ch6_A_wire\
        );

    \ch6_A_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39352\,
            PADOUT => \N__39351\,
            PADIN => \N__39350\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch6_A_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch6_B_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39343\,
            DIN => \N__39342\,
            DOUT => \N__39341\,
            PACKAGEPIN => \ch6_B_wire\
        );

    \ch6_B_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39343\,
            PADOUT => \N__39342\,
            PADIN => \N__39341\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch6_B_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch5_B_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39334\,
            DIN => \N__39333\,
            DOUT => \N__39332\,
            PACKAGEPIN => \ch5_B_wire\
        );

    \ch5_B_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39334\,
            PADOUT => \N__39333\,
            PADIN => \N__39332\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch5_B_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch0_B_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39325\,
            DIN => \N__39324\,
            DOUT => \N__39323\,
            PACKAGEPIN => \ch0_B_wire\
        );

    \ch0_B_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39325\,
            PADOUT => \N__39324\,
            PADIN => \N__39323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch0_B_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWM6_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39316\,
            DIN => \N__39315\,
            DOUT => \N__39314\,
            PACKAGEPIN => \PWM6_wire\
        );

    \PWM6_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39316\,
            PADOUT => \N__39315\,
            PADIN => \N__39314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__17397\,
            DIN0 => OPEN,
            DOUT0 => \N__21378\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWM4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39307\,
            DIN => \N__39306\,
            DOUT => \N__39305\,
            PACKAGEPIN => \PWM4_wire\
        );

    \PWM4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39307\,
            PADOUT => \N__39306\,
            PADIN => \N__39305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__27090\,
            DIN0 => OPEN,
            DOUT0 => \N__24981\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39298\,
            DIN => \N__39297\,
            DOUT => \N__39296\,
            PACKAGEPIN => \RST_wire\
        );

    \RST_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39298\,
            PADOUT => \N__39297\,
            PADIN => \N__39296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MISO_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39289\,
            DIN => \N__39288\,
            DOUT => \N__39287\,
            PACKAGEPIN => \MISO_wire\
        );

    \MISO_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39289\,
            PADOUT => \N__39288\,
            PADIN => \N__39287\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__36942\,
            DIN0 => OPEN,
            DOUT0 => \N__36639\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch5_A_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39280\,
            DIN => \N__39279\,
            DOUT => \N__39278\,
            PACKAGEPIN => \ch5_A_wire\
        );

    \ch5_A_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39280\,
            PADOUT => \N__39279\,
            PADIN => \N__39278\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch5_A_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch2_B_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39271\,
            DIN => \N__39270\,
            DOUT => \N__39269\,
            PACKAGEPIN => \ch2_B_wire\
        );

    \ch2_B_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39271\,
            PADOUT => \N__39270\,
            PADIN => \N__39269\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch2_B_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch4_B_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39262\,
            DIN => \N__39261\,
            DOUT => \N__39260\,
            PACKAGEPIN => \ch4_B_wire\
        );

    \ch4_B_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39262\,
            PADOUT => \N__39261\,
            PADIN => \N__39260\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch4_B_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWM3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39253\,
            DIN => \N__39252\,
            DOUT => \N__39251\,
            PACKAGEPIN => \PWM3_wire\
        );

    \PWM3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39253\,
            PADOUT => \N__39252\,
            PADIN => \N__39251\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__36948\,
            DIN0 => OPEN,
            DOUT0 => \N__29727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWM1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39244\,
            DIN => \N__39243\,
            DOUT => \N__39242\,
            PACKAGEPIN => \PWM1_wire\
        );

    \PWM1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39244\,
            PADOUT => \N__39243\,
            PADIN => \N__39242\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__17403\,
            DIN0 => OPEN,
            DOUT0 => \N__15735\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch4_A_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39235\,
            DIN => \N__39234\,
            DOUT => \N__39233\,
            PACKAGEPIN => \ch4_A_wire\
        );

    \ch4_A_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39235\,
            PADOUT => \N__39234\,
            PADIN => \N__39233\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch4_A_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch7_A_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39226\,
            DIN => \N__39225\,
            DOUT => \N__39224\,
            PACKAGEPIN => \ch7_A_wire\
        );

    \ch7_A_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39226\,
            PADOUT => \N__39225\,
            PADIN => \N__39224\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch7_A_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch3_B_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39217\,
            DIN => \N__39216\,
            DOUT => \N__39215\,
            PACKAGEPIN => \ch3_B_wire\
        );

    \ch3_B_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39217\,
            PADOUT => \N__39216\,
            PADIN => \N__39215\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch3_B_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWM7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39208\,
            DIN => \N__39207\,
            DOUT => \N__39206\,
            PACKAGEPIN => \PWM7_wire\
        );

    \PWM7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39208\,
            PADOUT => \N__39207\,
            PADIN => \N__39206\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__17391\,
            DIN0 => OPEN,
            DOUT0 => \N__14895\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39199\,
            DIN => \N__39198\,
            DOUT => \N__39197\,
            PACKAGEPIN => \SCK_wire\
        );

    \SCK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39199\,
            PADOUT => \N__39198\,
            PADIN => \N__39197\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SCK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch3_A_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39190\,
            DIN => \N__39189\,
            DOUT => \N__39188\,
            PACKAGEPIN => \ch3_A_wire\
        );

    \ch3_A_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39190\,
            PADOUT => \N__39189\,
            PADIN => \N__39188\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch3_A_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch1_B_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39181\,
            DIN => \N__39180\,
            DOUT => \N__39179\,
            PACKAGEPIN => \ch1_B_wire\
        );

    \ch1_B_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39181\,
            PADOUT => \N__39180\,
            PADIN => \N__39179\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch1_B_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWM2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39172\,
            DIN => \N__39171\,
            DOUT => \N__39170\,
            PACKAGEPIN => \PWM2_wire\
        );

    \PWM2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39172\,
            PADOUT => \N__39171\,
            PADIN => \N__39170\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35463\,
            DIN0 => OPEN,
            DOUT0 => \N__32151\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MOSI_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39163\,
            DIN => \N__39162\,
            DOUT => \N__39161\,
            PACKAGEPIN => \MOSI_wire\
        );

    \MOSI_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39163\,
            PADOUT => \N__39162\,
            PADIN => \N__39161\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \MOSI_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch7_B_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39154\,
            DIN => \N__39153\,
            DOUT => \N__39152\,
            PACKAGEPIN => \ch7_B_wire\
        );

    \ch7_B_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39154\,
            PADOUT => \N__39153\,
            PADIN => \N__39152\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch7_B_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch0_A_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39145\,
            DIN => \N__39144\,
            DOUT => \N__39143\,
            PACKAGEPIN => \ch0_A_wire\
        );

    \ch0_A_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39145\,
            PADOUT => \N__39144\,
            PADIN => \N__39143\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch0_A_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWM0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39136\,
            DIN => \N__39135\,
            DOUT => \N__39134\,
            PACKAGEPIN => \PWM0_wire\
        );

    \PWM0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39136\,
            PADOUT => \N__39135\,
            PADIN => \N__39134\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__17409\,
            DIN0 => OPEN,
            DOUT0 => \N__17250\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SSEL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39127\,
            DIN => \N__39126\,
            DOUT => \N__39125\,
            PACKAGEPIN => \SSEL_wire\
        );

    \SSEL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39127\,
            PADOUT => \N__39126\,
            PADIN => \N__39125\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SSEL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch1_A_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39118\,
            DIN => \N__39117\,
            DOUT => \N__39116\,
            PACKAGEPIN => \ch1_A_wire\
        );

    \ch1_A_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39118\,
            PADOUT => \N__39117\,
            PADIN => \N__39116\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch1_A_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ch2_A_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39109\,
            DIN => \N__39108\,
            DOUT => \N__39107\,
            PACKAGEPIN => \ch2_A_wire\
        );

    \ch2_A_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39109\,
            PADOUT => \N__39108\,
            PADIN => \N__39107\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ch2_A_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__9448\ : CascadeMux
    port map (
            O => \N__39090\,
            I => \N__39087\
        );

    \I__9447\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39084\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__39084\,
            I => \bit_count_RNIU615_0Z0Z_4\
        );

    \I__9445\ : CascadeMux
    port map (
            O => \N__39081\,
            I => \bit_count_RNIU615_0Z0Z_4_cascade_\
        );

    \I__9444\ : InMux
    port map (
            O => \N__39078\,
            I => \N__39075\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__39075\,
            I => \N__39072\
        );

    \I__9442\ : Span4Mux_h
    port map (
            O => \N__39072\,
            I => \N__39069\
        );

    \I__9441\ : Odrv4
    port map (
            O => \N__39069\,
            I => \SSELr_RNIGO0FZ0Z_1\
        );

    \I__9440\ : InMux
    port map (
            O => \N__39066\,
            I => \N__39057\
        );

    \I__9439\ : InMux
    port map (
            O => \N__39065\,
            I => \N__39057\
        );

    \I__9438\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39057\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__39057\,
            I => \N__39050\
        );

    \I__9436\ : InMux
    port map (
            O => \N__39056\,
            I => \N__39037\
        );

    \I__9435\ : InMux
    port map (
            O => \N__39055\,
            I => \N__39037\
        );

    \I__9434\ : InMux
    port map (
            O => \N__39054\,
            I => \N__39037\
        );

    \I__9433\ : InMux
    port map (
            O => \N__39053\,
            I => \N__39037\
        );

    \I__9432\ : Span4Mux_h
    port map (
            O => \N__39050\,
            I => \N__39031\
        );

    \I__9431\ : InMux
    port map (
            O => \N__39049\,
            I => \N__39024\
        );

    \I__9430\ : InMux
    port map (
            O => \N__39048\,
            I => \N__39024\
        );

    \I__9429\ : InMux
    port map (
            O => \N__39047\,
            I => \N__39024\
        );

    \I__9428\ : InMux
    port map (
            O => \N__39046\,
            I => \N__39021\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__39037\,
            I => \N__39018\
        );

    \I__9426\ : InMux
    port map (
            O => \N__39036\,
            I => \N__39011\
        );

    \I__9425\ : InMux
    port map (
            O => \N__39035\,
            I => \N__39011\
        );

    \I__9424\ : InMux
    port map (
            O => \N__39034\,
            I => \N__39011\
        );

    \I__9423\ : Span4Mux_h
    port map (
            O => \N__39031\,
            I => \N__39006\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__39024\,
            I => \N__39006\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__39021\,
            I => \SSELrZ0Z_1\
        );

    \I__9420\ : Odrv12
    port map (
            O => \N__39018\,
            I => \SSELrZ0Z_1\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__39011\,
            I => \SSELrZ0Z_1\
        );

    \I__9418\ : Odrv4
    port map (
            O => \N__39006\,
            I => \SSELrZ0Z_1\
        );

    \I__9417\ : CascadeMux
    port map (
            O => \N__38997\,
            I => \N__38994\
        );

    \I__9416\ : InMux
    port map (
            O => \N__38994\,
            I => \N__38988\
        );

    \I__9415\ : InMux
    port map (
            O => \N__38993\,
            I => \N__38988\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__38988\,
            I => un1_bit_count_1_c3
        );

    \I__9413\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38979\
        );

    \I__9412\ : InMux
    port map (
            O => \N__38984\,
            I => \N__38972\
        );

    \I__9411\ : InMux
    port map (
            O => \N__38983\,
            I => \N__38972\
        );

    \I__9410\ : InMux
    port map (
            O => \N__38982\,
            I => \N__38972\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__38979\,
            I => \bit_countZ0Z_3\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__38972\,
            I => \bit_countZ0Z_3\
        );

    \I__9407\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38962\
        );

    \I__9406\ : InMux
    port map (
            O => \N__38966\,
            I => \N__38957\
        );

    \I__9405\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38957\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__38962\,
            I => \bit_countZ0Z_4\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__38957\,
            I => \bit_countZ0Z_4\
        );

    \I__9402\ : CascadeMux
    port map (
            O => \N__38952\,
            I => \N__38948\
        );

    \I__9401\ : InMux
    port map (
            O => \N__38951\,
            I => \N__38943\
        );

    \I__9400\ : InMux
    port map (
            O => \N__38948\,
            I => \N__38938\
        );

    \I__9399\ : InMux
    port map (
            O => \N__38947\,
            I => \N__38938\
        );

    \I__9398\ : InMux
    port map (
            O => \N__38946\,
            I => \N__38934\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__38943\,
            I => \N__38929\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__38938\,
            I => \N__38926\
        );

    \I__9395\ : InMux
    port map (
            O => \N__38937\,
            I => \N__38923\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__38934\,
            I => \N__38920\
        );

    \I__9393\ : InMux
    port map (
            O => \N__38933\,
            I => \N__38917\
        );

    \I__9392\ : InMux
    port map (
            O => \N__38932\,
            I => \N__38914\
        );

    \I__9391\ : Span4Mux_v
    port map (
            O => \N__38929\,
            I => \N__38905\
        );

    \I__9390\ : Span4Mux_v
    port map (
            O => \N__38926\,
            I => \N__38905\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__38923\,
            I => \N__38902\
        );

    \I__9388\ : Span4Mux_h
    port map (
            O => \N__38920\,
            I => \N__38893\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__38917\,
            I => \N__38893\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__38914\,
            I => \N__38893\
        );

    \I__9385\ : InMux
    port map (
            O => \N__38913\,
            I => \N__38890\
        );

    \I__9384\ : InMux
    port map (
            O => \N__38912\,
            I => \N__38887\
        );

    \I__9383\ : CascadeMux
    port map (
            O => \N__38911\,
            I => \N__38884\
        );

    \I__9382\ : CascadeMux
    port map (
            O => \N__38910\,
            I => \N__38880\
        );

    \I__9381\ : Span4Mux_h
    port map (
            O => \N__38905\,
            I => \N__38872\
        );

    \I__9380\ : Span4Mux_h
    port map (
            O => \N__38902\,
            I => \N__38872\
        );

    \I__9379\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38869\
        );

    \I__9378\ : InMux
    port map (
            O => \N__38900\,
            I => \N__38866\
        );

    \I__9377\ : Span4Mux_v
    port map (
            O => \N__38893\,
            I => \N__38857\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__38890\,
            I => \N__38857\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__38887\,
            I => \N__38857\
        );

    \I__9374\ : InMux
    port map (
            O => \N__38884\,
            I => \N__38852\
        );

    \I__9373\ : InMux
    port map (
            O => \N__38883\,
            I => \N__38852\
        );

    \I__9372\ : InMux
    port map (
            O => \N__38880\,
            I => \N__38847\
        );

    \I__9371\ : InMux
    port map (
            O => \N__38879\,
            I => \N__38847\
        );

    \I__9370\ : InMux
    port map (
            O => \N__38878\,
            I => \N__38842\
        );

    \I__9369\ : InMux
    port map (
            O => \N__38877\,
            I => \N__38842\
        );

    \I__9368\ : Span4Mux_h
    port map (
            O => \N__38872\,
            I => \N__38837\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__38869\,
            I => \N__38837\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__38866\,
            I => \N__38834\
        );

    \I__9365\ : InMux
    port map (
            O => \N__38865\,
            I => \N__38831\
        );

    \I__9364\ : InMux
    port map (
            O => \N__38864\,
            I => \N__38828\
        );

    \I__9363\ : Span4Mux_h
    port map (
            O => \N__38857\,
            I => \N__38825\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__38852\,
            I => \N__38818\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__38847\,
            I => \N__38818\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__38842\,
            I => \N__38818\
        );

    \I__9359\ : Odrv4
    port map (
            O => \N__38837\,
            I => \un1_OutReg51_4_0_i_o3_3\
        );

    \I__9358\ : Odrv4
    port map (
            O => \N__38834\,
            I => \un1_OutReg51_4_0_i_o3_3\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__38831\,
            I => \un1_OutReg51_4_0_i_o3_3\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__38828\,
            I => \un1_OutReg51_4_0_i_o3_3\
        );

    \I__9355\ : Odrv4
    port map (
            O => \N__38825\,
            I => \un1_OutReg51_4_0_i_o3_3\
        );

    \I__9354\ : Odrv12
    port map (
            O => \N__38818\,
            I => \un1_OutReg51_4_0_i_o3_3\
        );

    \I__9353\ : CascadeMux
    port map (
            O => \N__38805\,
            I => \N__38802\
        );

    \I__9352\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38799\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__38799\,
            I => \N__38790\
        );

    \I__9350\ : InMux
    port map (
            O => \N__38798\,
            I => \N__38787\
        );

    \I__9349\ : InMux
    port map (
            O => \N__38797\,
            I => \N__38782\
        );

    \I__9348\ : InMux
    port map (
            O => \N__38796\,
            I => \N__38782\
        );

    \I__9347\ : InMux
    port map (
            O => \N__38795\,
            I => \N__38777\
        );

    \I__9346\ : InMux
    port map (
            O => \N__38794\,
            I => \N__38777\
        );

    \I__9345\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38774\
        );

    \I__9344\ : Odrv4
    port map (
            O => \N__38790\,
            I => \SCKrZ0Z_1\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__38787\,
            I => \SCKrZ0Z_1\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__38782\,
            I => \SCKrZ0Z_1\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__38777\,
            I => \SCKrZ0Z_1\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__38774\,
            I => \SCKrZ0Z_1\
        );

    \I__9339\ : CascadeMux
    port map (
            O => \N__38763\,
            I => \N__38755\
        );

    \I__9338\ : CascadeMux
    port map (
            O => \N__38762\,
            I => \N__38752\
        );

    \I__9337\ : InMux
    port map (
            O => \N__38761\,
            I => \N__38747\
        );

    \I__9336\ : InMux
    port map (
            O => \N__38760\,
            I => \N__38747\
        );

    \I__9335\ : InMux
    port map (
            O => \N__38759\,
            I => \N__38744\
        );

    \I__9334\ : InMux
    port map (
            O => \N__38758\,
            I => \N__38741\
        );

    \I__9333\ : InMux
    port map (
            O => \N__38755\,
            I => \N__38738\
        );

    \I__9332\ : InMux
    port map (
            O => \N__38752\,
            I => \N__38735\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__38747\,
            I => \SCKrZ0Z_2\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__38744\,
            I => \SCKrZ0Z_2\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__38741\,
            I => \SCKrZ0Z_2\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__38738\,
            I => \SCKrZ0Z_2\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__38735\,
            I => \SCKrZ0Z_2\
        );

    \I__9326\ : ClkMux
    port map (
            O => \N__38724\,
            I => \N__38172\
        );

    \I__9325\ : ClkMux
    port map (
            O => \N__38723\,
            I => \N__38172\
        );

    \I__9324\ : ClkMux
    port map (
            O => \N__38722\,
            I => \N__38172\
        );

    \I__9323\ : ClkMux
    port map (
            O => \N__38721\,
            I => \N__38172\
        );

    \I__9322\ : ClkMux
    port map (
            O => \N__38720\,
            I => \N__38172\
        );

    \I__9321\ : ClkMux
    port map (
            O => \N__38719\,
            I => \N__38172\
        );

    \I__9320\ : ClkMux
    port map (
            O => \N__38718\,
            I => \N__38172\
        );

    \I__9319\ : ClkMux
    port map (
            O => \N__38717\,
            I => \N__38172\
        );

    \I__9318\ : ClkMux
    port map (
            O => \N__38716\,
            I => \N__38172\
        );

    \I__9317\ : ClkMux
    port map (
            O => \N__38715\,
            I => \N__38172\
        );

    \I__9316\ : ClkMux
    port map (
            O => \N__38714\,
            I => \N__38172\
        );

    \I__9315\ : ClkMux
    port map (
            O => \N__38713\,
            I => \N__38172\
        );

    \I__9314\ : ClkMux
    port map (
            O => \N__38712\,
            I => \N__38172\
        );

    \I__9313\ : ClkMux
    port map (
            O => \N__38711\,
            I => \N__38172\
        );

    \I__9312\ : ClkMux
    port map (
            O => \N__38710\,
            I => \N__38172\
        );

    \I__9311\ : ClkMux
    port map (
            O => \N__38709\,
            I => \N__38172\
        );

    \I__9310\ : ClkMux
    port map (
            O => \N__38708\,
            I => \N__38172\
        );

    \I__9309\ : ClkMux
    port map (
            O => \N__38707\,
            I => \N__38172\
        );

    \I__9308\ : ClkMux
    port map (
            O => \N__38706\,
            I => \N__38172\
        );

    \I__9307\ : ClkMux
    port map (
            O => \N__38705\,
            I => \N__38172\
        );

    \I__9306\ : ClkMux
    port map (
            O => \N__38704\,
            I => \N__38172\
        );

    \I__9305\ : ClkMux
    port map (
            O => \N__38703\,
            I => \N__38172\
        );

    \I__9304\ : ClkMux
    port map (
            O => \N__38702\,
            I => \N__38172\
        );

    \I__9303\ : ClkMux
    port map (
            O => \N__38701\,
            I => \N__38172\
        );

    \I__9302\ : ClkMux
    port map (
            O => \N__38700\,
            I => \N__38172\
        );

    \I__9301\ : ClkMux
    port map (
            O => \N__38699\,
            I => \N__38172\
        );

    \I__9300\ : ClkMux
    port map (
            O => \N__38698\,
            I => \N__38172\
        );

    \I__9299\ : ClkMux
    port map (
            O => \N__38697\,
            I => \N__38172\
        );

    \I__9298\ : ClkMux
    port map (
            O => \N__38696\,
            I => \N__38172\
        );

    \I__9297\ : ClkMux
    port map (
            O => \N__38695\,
            I => \N__38172\
        );

    \I__9296\ : ClkMux
    port map (
            O => \N__38694\,
            I => \N__38172\
        );

    \I__9295\ : ClkMux
    port map (
            O => \N__38693\,
            I => \N__38172\
        );

    \I__9294\ : ClkMux
    port map (
            O => \N__38692\,
            I => \N__38172\
        );

    \I__9293\ : ClkMux
    port map (
            O => \N__38691\,
            I => \N__38172\
        );

    \I__9292\ : ClkMux
    port map (
            O => \N__38690\,
            I => \N__38172\
        );

    \I__9291\ : ClkMux
    port map (
            O => \N__38689\,
            I => \N__38172\
        );

    \I__9290\ : ClkMux
    port map (
            O => \N__38688\,
            I => \N__38172\
        );

    \I__9289\ : ClkMux
    port map (
            O => \N__38687\,
            I => \N__38172\
        );

    \I__9288\ : ClkMux
    port map (
            O => \N__38686\,
            I => \N__38172\
        );

    \I__9287\ : ClkMux
    port map (
            O => \N__38685\,
            I => \N__38172\
        );

    \I__9286\ : ClkMux
    port map (
            O => \N__38684\,
            I => \N__38172\
        );

    \I__9285\ : ClkMux
    port map (
            O => \N__38683\,
            I => \N__38172\
        );

    \I__9284\ : ClkMux
    port map (
            O => \N__38682\,
            I => \N__38172\
        );

    \I__9283\ : ClkMux
    port map (
            O => \N__38681\,
            I => \N__38172\
        );

    \I__9282\ : ClkMux
    port map (
            O => \N__38680\,
            I => \N__38172\
        );

    \I__9281\ : ClkMux
    port map (
            O => \N__38679\,
            I => \N__38172\
        );

    \I__9280\ : ClkMux
    port map (
            O => \N__38678\,
            I => \N__38172\
        );

    \I__9279\ : ClkMux
    port map (
            O => \N__38677\,
            I => \N__38172\
        );

    \I__9278\ : ClkMux
    port map (
            O => \N__38676\,
            I => \N__38172\
        );

    \I__9277\ : ClkMux
    port map (
            O => \N__38675\,
            I => \N__38172\
        );

    \I__9276\ : ClkMux
    port map (
            O => \N__38674\,
            I => \N__38172\
        );

    \I__9275\ : ClkMux
    port map (
            O => \N__38673\,
            I => \N__38172\
        );

    \I__9274\ : ClkMux
    port map (
            O => \N__38672\,
            I => \N__38172\
        );

    \I__9273\ : ClkMux
    port map (
            O => \N__38671\,
            I => \N__38172\
        );

    \I__9272\ : ClkMux
    port map (
            O => \N__38670\,
            I => \N__38172\
        );

    \I__9271\ : ClkMux
    port map (
            O => \N__38669\,
            I => \N__38172\
        );

    \I__9270\ : ClkMux
    port map (
            O => \N__38668\,
            I => \N__38172\
        );

    \I__9269\ : ClkMux
    port map (
            O => \N__38667\,
            I => \N__38172\
        );

    \I__9268\ : ClkMux
    port map (
            O => \N__38666\,
            I => \N__38172\
        );

    \I__9267\ : ClkMux
    port map (
            O => \N__38665\,
            I => \N__38172\
        );

    \I__9266\ : ClkMux
    port map (
            O => \N__38664\,
            I => \N__38172\
        );

    \I__9265\ : ClkMux
    port map (
            O => \N__38663\,
            I => \N__38172\
        );

    \I__9264\ : ClkMux
    port map (
            O => \N__38662\,
            I => \N__38172\
        );

    \I__9263\ : ClkMux
    port map (
            O => \N__38661\,
            I => \N__38172\
        );

    \I__9262\ : ClkMux
    port map (
            O => \N__38660\,
            I => \N__38172\
        );

    \I__9261\ : ClkMux
    port map (
            O => \N__38659\,
            I => \N__38172\
        );

    \I__9260\ : ClkMux
    port map (
            O => \N__38658\,
            I => \N__38172\
        );

    \I__9259\ : ClkMux
    port map (
            O => \N__38657\,
            I => \N__38172\
        );

    \I__9258\ : ClkMux
    port map (
            O => \N__38656\,
            I => \N__38172\
        );

    \I__9257\ : ClkMux
    port map (
            O => \N__38655\,
            I => \N__38172\
        );

    \I__9256\ : ClkMux
    port map (
            O => \N__38654\,
            I => \N__38172\
        );

    \I__9255\ : ClkMux
    port map (
            O => \N__38653\,
            I => \N__38172\
        );

    \I__9254\ : ClkMux
    port map (
            O => \N__38652\,
            I => \N__38172\
        );

    \I__9253\ : ClkMux
    port map (
            O => \N__38651\,
            I => \N__38172\
        );

    \I__9252\ : ClkMux
    port map (
            O => \N__38650\,
            I => \N__38172\
        );

    \I__9251\ : ClkMux
    port map (
            O => \N__38649\,
            I => \N__38172\
        );

    \I__9250\ : ClkMux
    port map (
            O => \N__38648\,
            I => \N__38172\
        );

    \I__9249\ : ClkMux
    port map (
            O => \N__38647\,
            I => \N__38172\
        );

    \I__9248\ : ClkMux
    port map (
            O => \N__38646\,
            I => \N__38172\
        );

    \I__9247\ : ClkMux
    port map (
            O => \N__38645\,
            I => \N__38172\
        );

    \I__9246\ : ClkMux
    port map (
            O => \N__38644\,
            I => \N__38172\
        );

    \I__9245\ : ClkMux
    port map (
            O => \N__38643\,
            I => \N__38172\
        );

    \I__9244\ : ClkMux
    port map (
            O => \N__38642\,
            I => \N__38172\
        );

    \I__9243\ : ClkMux
    port map (
            O => \N__38641\,
            I => \N__38172\
        );

    \I__9242\ : ClkMux
    port map (
            O => \N__38640\,
            I => \N__38172\
        );

    \I__9241\ : ClkMux
    port map (
            O => \N__38639\,
            I => \N__38172\
        );

    \I__9240\ : ClkMux
    port map (
            O => \N__38638\,
            I => \N__38172\
        );

    \I__9239\ : ClkMux
    port map (
            O => \N__38637\,
            I => \N__38172\
        );

    \I__9238\ : ClkMux
    port map (
            O => \N__38636\,
            I => \N__38172\
        );

    \I__9237\ : ClkMux
    port map (
            O => \N__38635\,
            I => \N__38172\
        );

    \I__9236\ : ClkMux
    port map (
            O => \N__38634\,
            I => \N__38172\
        );

    \I__9235\ : ClkMux
    port map (
            O => \N__38633\,
            I => \N__38172\
        );

    \I__9234\ : ClkMux
    port map (
            O => \N__38632\,
            I => \N__38172\
        );

    \I__9233\ : ClkMux
    port map (
            O => \N__38631\,
            I => \N__38172\
        );

    \I__9232\ : ClkMux
    port map (
            O => \N__38630\,
            I => \N__38172\
        );

    \I__9231\ : ClkMux
    port map (
            O => \N__38629\,
            I => \N__38172\
        );

    \I__9230\ : ClkMux
    port map (
            O => \N__38628\,
            I => \N__38172\
        );

    \I__9229\ : ClkMux
    port map (
            O => \N__38627\,
            I => \N__38172\
        );

    \I__9228\ : ClkMux
    port map (
            O => \N__38626\,
            I => \N__38172\
        );

    \I__9227\ : ClkMux
    port map (
            O => \N__38625\,
            I => \N__38172\
        );

    \I__9226\ : ClkMux
    port map (
            O => \N__38624\,
            I => \N__38172\
        );

    \I__9225\ : ClkMux
    port map (
            O => \N__38623\,
            I => \N__38172\
        );

    \I__9224\ : ClkMux
    port map (
            O => \N__38622\,
            I => \N__38172\
        );

    \I__9223\ : ClkMux
    port map (
            O => \N__38621\,
            I => \N__38172\
        );

    \I__9222\ : ClkMux
    port map (
            O => \N__38620\,
            I => \N__38172\
        );

    \I__9221\ : ClkMux
    port map (
            O => \N__38619\,
            I => \N__38172\
        );

    \I__9220\ : ClkMux
    port map (
            O => \N__38618\,
            I => \N__38172\
        );

    \I__9219\ : ClkMux
    port map (
            O => \N__38617\,
            I => \N__38172\
        );

    \I__9218\ : ClkMux
    port map (
            O => \N__38616\,
            I => \N__38172\
        );

    \I__9217\ : ClkMux
    port map (
            O => \N__38615\,
            I => \N__38172\
        );

    \I__9216\ : ClkMux
    port map (
            O => \N__38614\,
            I => \N__38172\
        );

    \I__9215\ : ClkMux
    port map (
            O => \N__38613\,
            I => \N__38172\
        );

    \I__9214\ : ClkMux
    port map (
            O => \N__38612\,
            I => \N__38172\
        );

    \I__9213\ : ClkMux
    port map (
            O => \N__38611\,
            I => \N__38172\
        );

    \I__9212\ : ClkMux
    port map (
            O => \N__38610\,
            I => \N__38172\
        );

    \I__9211\ : ClkMux
    port map (
            O => \N__38609\,
            I => \N__38172\
        );

    \I__9210\ : ClkMux
    port map (
            O => \N__38608\,
            I => \N__38172\
        );

    \I__9209\ : ClkMux
    port map (
            O => \N__38607\,
            I => \N__38172\
        );

    \I__9208\ : ClkMux
    port map (
            O => \N__38606\,
            I => \N__38172\
        );

    \I__9207\ : ClkMux
    port map (
            O => \N__38605\,
            I => \N__38172\
        );

    \I__9206\ : ClkMux
    port map (
            O => \N__38604\,
            I => \N__38172\
        );

    \I__9205\ : ClkMux
    port map (
            O => \N__38603\,
            I => \N__38172\
        );

    \I__9204\ : ClkMux
    port map (
            O => \N__38602\,
            I => \N__38172\
        );

    \I__9203\ : ClkMux
    port map (
            O => \N__38601\,
            I => \N__38172\
        );

    \I__9202\ : ClkMux
    port map (
            O => \N__38600\,
            I => \N__38172\
        );

    \I__9201\ : ClkMux
    port map (
            O => \N__38599\,
            I => \N__38172\
        );

    \I__9200\ : ClkMux
    port map (
            O => \N__38598\,
            I => \N__38172\
        );

    \I__9199\ : ClkMux
    port map (
            O => \N__38597\,
            I => \N__38172\
        );

    \I__9198\ : ClkMux
    port map (
            O => \N__38596\,
            I => \N__38172\
        );

    \I__9197\ : ClkMux
    port map (
            O => \N__38595\,
            I => \N__38172\
        );

    \I__9196\ : ClkMux
    port map (
            O => \N__38594\,
            I => \N__38172\
        );

    \I__9195\ : ClkMux
    port map (
            O => \N__38593\,
            I => \N__38172\
        );

    \I__9194\ : ClkMux
    port map (
            O => \N__38592\,
            I => \N__38172\
        );

    \I__9193\ : ClkMux
    port map (
            O => \N__38591\,
            I => \N__38172\
        );

    \I__9192\ : ClkMux
    port map (
            O => \N__38590\,
            I => \N__38172\
        );

    \I__9191\ : ClkMux
    port map (
            O => \N__38589\,
            I => \N__38172\
        );

    \I__9190\ : ClkMux
    port map (
            O => \N__38588\,
            I => \N__38172\
        );

    \I__9189\ : ClkMux
    port map (
            O => \N__38587\,
            I => \N__38172\
        );

    \I__9188\ : ClkMux
    port map (
            O => \N__38586\,
            I => \N__38172\
        );

    \I__9187\ : ClkMux
    port map (
            O => \N__38585\,
            I => \N__38172\
        );

    \I__9186\ : ClkMux
    port map (
            O => \N__38584\,
            I => \N__38172\
        );

    \I__9185\ : ClkMux
    port map (
            O => \N__38583\,
            I => \N__38172\
        );

    \I__9184\ : ClkMux
    port map (
            O => \N__38582\,
            I => \N__38172\
        );

    \I__9183\ : ClkMux
    port map (
            O => \N__38581\,
            I => \N__38172\
        );

    \I__9182\ : ClkMux
    port map (
            O => \N__38580\,
            I => \N__38172\
        );

    \I__9181\ : ClkMux
    port map (
            O => \N__38579\,
            I => \N__38172\
        );

    \I__9180\ : ClkMux
    port map (
            O => \N__38578\,
            I => \N__38172\
        );

    \I__9179\ : ClkMux
    port map (
            O => \N__38577\,
            I => \N__38172\
        );

    \I__9178\ : ClkMux
    port map (
            O => \N__38576\,
            I => \N__38172\
        );

    \I__9177\ : ClkMux
    port map (
            O => \N__38575\,
            I => \N__38172\
        );

    \I__9176\ : ClkMux
    port map (
            O => \N__38574\,
            I => \N__38172\
        );

    \I__9175\ : ClkMux
    port map (
            O => \N__38573\,
            I => \N__38172\
        );

    \I__9174\ : ClkMux
    port map (
            O => \N__38572\,
            I => \N__38172\
        );

    \I__9173\ : ClkMux
    port map (
            O => \N__38571\,
            I => \N__38172\
        );

    \I__9172\ : ClkMux
    port map (
            O => \N__38570\,
            I => \N__38172\
        );

    \I__9171\ : ClkMux
    port map (
            O => \N__38569\,
            I => \N__38172\
        );

    \I__9170\ : ClkMux
    port map (
            O => \N__38568\,
            I => \N__38172\
        );

    \I__9169\ : ClkMux
    port map (
            O => \N__38567\,
            I => \N__38172\
        );

    \I__9168\ : ClkMux
    port map (
            O => \N__38566\,
            I => \N__38172\
        );

    \I__9167\ : ClkMux
    port map (
            O => \N__38565\,
            I => \N__38172\
        );

    \I__9166\ : ClkMux
    port map (
            O => \N__38564\,
            I => \N__38172\
        );

    \I__9165\ : ClkMux
    port map (
            O => \N__38563\,
            I => \N__38172\
        );

    \I__9164\ : ClkMux
    port map (
            O => \N__38562\,
            I => \N__38172\
        );

    \I__9163\ : ClkMux
    port map (
            O => \N__38561\,
            I => \N__38172\
        );

    \I__9162\ : ClkMux
    port map (
            O => \N__38560\,
            I => \N__38172\
        );

    \I__9161\ : ClkMux
    port map (
            O => \N__38559\,
            I => \N__38172\
        );

    \I__9160\ : ClkMux
    port map (
            O => \N__38558\,
            I => \N__38172\
        );

    \I__9159\ : ClkMux
    port map (
            O => \N__38557\,
            I => \N__38172\
        );

    \I__9158\ : ClkMux
    port map (
            O => \N__38556\,
            I => \N__38172\
        );

    \I__9157\ : ClkMux
    port map (
            O => \N__38555\,
            I => \N__38172\
        );

    \I__9156\ : ClkMux
    port map (
            O => \N__38554\,
            I => \N__38172\
        );

    \I__9155\ : ClkMux
    port map (
            O => \N__38553\,
            I => \N__38172\
        );

    \I__9154\ : ClkMux
    port map (
            O => \N__38552\,
            I => \N__38172\
        );

    \I__9153\ : ClkMux
    port map (
            O => \N__38551\,
            I => \N__38172\
        );

    \I__9152\ : ClkMux
    port map (
            O => \N__38550\,
            I => \N__38172\
        );

    \I__9151\ : ClkMux
    port map (
            O => \N__38549\,
            I => \N__38172\
        );

    \I__9150\ : ClkMux
    port map (
            O => \N__38548\,
            I => \N__38172\
        );

    \I__9149\ : ClkMux
    port map (
            O => \N__38547\,
            I => \N__38172\
        );

    \I__9148\ : ClkMux
    port map (
            O => \N__38546\,
            I => \N__38172\
        );

    \I__9147\ : ClkMux
    port map (
            O => \N__38545\,
            I => \N__38172\
        );

    \I__9146\ : ClkMux
    port map (
            O => \N__38544\,
            I => \N__38172\
        );

    \I__9145\ : ClkMux
    port map (
            O => \N__38543\,
            I => \N__38172\
        );

    \I__9144\ : ClkMux
    port map (
            O => \N__38542\,
            I => \N__38172\
        );

    \I__9143\ : ClkMux
    port map (
            O => \N__38541\,
            I => \N__38172\
        );

    \I__9142\ : GlobalMux
    port map (
            O => \N__38172\,
            I => \N__38169\
        );

    \I__9141\ : gio2CtrlBuf
    port map (
            O => \N__38169\,
            I => myclk
        );

    \I__9140\ : CascadeMux
    port map (
            O => \N__38166\,
            I => \N__38163\
        );

    \I__9139\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38160\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__38160\,
            I => \N__38149\
        );

    \I__9137\ : InMux
    port map (
            O => \N__38159\,
            I => \N__38146\
        );

    \I__9136\ : InMux
    port map (
            O => \N__38158\,
            I => \N__38143\
        );

    \I__9135\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38140\
        );

    \I__9134\ : InMux
    port map (
            O => \N__38156\,
            I => \N__38132\
        );

    \I__9133\ : InMux
    port map (
            O => \N__38155\,
            I => \N__38132\
        );

    \I__9132\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38129\
        );

    \I__9131\ : InMux
    port map (
            O => \N__38153\,
            I => \N__38126\
        );

    \I__9130\ : InMux
    port map (
            O => \N__38152\,
            I => \N__38123\
        );

    \I__9129\ : Span4Mux_h
    port map (
            O => \N__38149\,
            I => \N__38118\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__38146\,
            I => \N__38118\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__38143\,
            I => \N__38115\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__38140\,
            I => \N__38110\
        );

    \I__9125\ : InMux
    port map (
            O => \N__38139\,
            I => \N__38107\
        );

    \I__9124\ : InMux
    port map (
            O => \N__38138\,
            I => \N__38104\
        );

    \I__9123\ : CascadeMux
    port map (
            O => \N__38137\,
            I => \N__38101\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__38132\,
            I => \N__38097\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__38129\,
            I => \N__38091\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__38126\,
            I => \N__38088\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__38123\,
            I => \N__38085\
        );

    \I__9118\ : Span4Mux_v
    port map (
            O => \N__38118\,
            I => \N__38080\
        );

    \I__9117\ : Span4Mux_h
    port map (
            O => \N__38115\,
            I => \N__38080\
        );

    \I__9116\ : InMux
    port map (
            O => \N__38114\,
            I => \N__38077\
        );

    \I__9115\ : InMux
    port map (
            O => \N__38113\,
            I => \N__38074\
        );

    \I__9114\ : Span4Mux_v
    port map (
            O => \N__38110\,
            I => \N__38067\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__38107\,
            I => \N__38067\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__38104\,
            I => \N__38067\
        );

    \I__9111\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38064\
        );

    \I__9110\ : InMux
    port map (
            O => \N__38100\,
            I => \N__38061\
        );

    \I__9109\ : Span4Mux_h
    port map (
            O => \N__38097\,
            I => \N__38058\
        );

    \I__9108\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38055\
        );

    \I__9107\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38052\
        );

    \I__9106\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38049\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__38091\,
            I => \N__38042\
        );

    \I__9104\ : Span4Mux_h
    port map (
            O => \N__38088\,
            I => \N__38042\
        );

    \I__9103\ : Span4Mux_h
    port map (
            O => \N__38085\,
            I => \N__38042\
        );

    \I__9102\ : Span4Mux_h
    port map (
            O => \N__38080\,
            I => \N__38037\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__38077\,
            I => \N__38037\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__38074\,
            I => \N__38030\
        );

    \I__9099\ : Span4Mux_h
    port map (
            O => \N__38067\,
            I => \N__38030\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__38064\,
            I => \N__38030\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__38061\,
            I => \data_receivedZ0Z_0\
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__38058\,
            I => \data_receivedZ0Z_0\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__38055\,
            I => \data_receivedZ0Z_0\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__38052\,
            I => \data_receivedZ0Z_0\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__38049\,
            I => \data_receivedZ0Z_0\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__38042\,
            I => \data_receivedZ0Z_0\
        );

    \I__9091\ : Odrv4
    port map (
            O => \N__38037\,
            I => \data_receivedZ0Z_0\
        );

    \I__9090\ : Odrv4
    port map (
            O => \N__38030\,
            I => \data_receivedZ0Z_0\
        );

    \I__9089\ : InMux
    port map (
            O => \N__38013\,
            I => \N__38010\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__38010\,
            I => \N__38007\
        );

    \I__9087\ : Span4Mux_v
    port map (
            O => \N__38007\,
            I => \N__38004\
        );

    \I__9086\ : Odrv4
    port map (
            O => \N__38004\,
            I => \OutReg_0_5_i_m3_ns_1_8\
        );

    \I__9085\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37998\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__37998\,
            I => \OutReg_esr_RNO_2Z0Z_8\
        );

    \I__9083\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37992\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__37992\,
            I => \N__37989\
        );

    \I__9081\ : Odrv4
    port map (
            O => \N__37989\,
            I => \SSELrZ0Z_0\
        );

    \I__9080\ : InMux
    port map (
            O => \N__37986\,
            I => \N__37977\
        );

    \I__9079\ : InMux
    port map (
            O => \N__37985\,
            I => \N__37977\
        );

    \I__9078\ : InMux
    port map (
            O => \N__37984\,
            I => \N__37977\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__37977\,
            I => \N__37974\
        );

    \I__9076\ : Odrv12
    port map (
            O => \N__37974\,
            I => \SSELrZ0Z_2\
        );

    \I__9075\ : InMux
    port map (
            O => \N__37971\,
            I => \N__37968\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__37968\,
            I => \N__37965\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__37965\,
            I => \SCK_c\
        );

    \I__9072\ : InMux
    port map (
            O => \N__37962\,
            I => \N__37957\
        );

    \I__9071\ : InMux
    port map (
            O => \N__37961\,
            I => \N__37954\
        );

    \I__9070\ : InMux
    port map (
            O => \N__37960\,
            I => \N__37951\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__37957\,
            I => \N__37946\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__37954\,
            I => \N__37946\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__37951\,
            I => \bit_countZ0Z_2\
        );

    \I__9066\ : Odrv4
    port map (
            O => \N__37946\,
            I => \bit_countZ0Z_2\
        );

    \I__9065\ : IoInMux
    port map (
            O => \N__37941\,
            I => \N__37938\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__37938\,
            I => \N__37935\
        );

    \I__9063\ : IoSpan4Mux
    port map (
            O => \N__37935\,
            I => \N__37932\
        );

    \I__9062\ : Sp12to4
    port map (
            O => \N__37932\,
            I => \N__37929\
        );

    \I__9061\ : Odrv12
    port map (
            O => \N__37929\,
            I => \SCKr_RNIBA7CZ0Z_2\
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__37926\,
            I => \SCKr_RNIBA7CZ0Z_2_cascade_\
        );

    \I__9059\ : IoInMux
    port map (
            O => \N__37923\,
            I => \N__37920\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__37920\,
            I => \N__37917\
        );

    \I__9057\ : Span4Mux_s0_v
    port map (
            O => \N__37917\,
            I => \N__37914\
        );

    \I__9056\ : Sp12to4
    port map (
            O => \N__37914\,
            I => \N__37911\
        );

    \I__9055\ : Span12Mux_h
    port map (
            O => \N__37911\,
            I => \N__37908\
        );

    \I__9054\ : Odrv12
    port map (
            O => \N__37908\,
            I => \N_45_0\
        );

    \I__9053\ : InMux
    port map (
            O => \N__37905\,
            I => \N__37902\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__37902\,
            I => \N__37899\
        );

    \I__9051\ : Odrv12
    port map (
            O => \N__37899\,
            I => \SCKrZ0Z_0\
        );

    \I__9050\ : InMux
    port map (
            O => \N__37896\,
            I => \N__37890\
        );

    \I__9049\ : InMux
    port map (
            O => \N__37895\,
            I => \N__37890\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__37890\,
            I => un1_bit_count_1_c1
        );

    \I__9047\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37881\
        );

    \I__9046\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37878\
        );

    \I__9045\ : InMux
    port map (
            O => \N__37885\,
            I => \N__37873\
        );

    \I__9044\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37873\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__37881\,
            I => \N__37868\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__37878\,
            I => \N__37868\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__37873\,
            I => \bit_countZ0Z_1\
        );

    \I__9040\ : Odrv4
    port map (
            O => \N__37868\,
            I => \bit_countZ0Z_1\
        );

    \I__9039\ : InMux
    port map (
            O => \N__37863\,
            I => \N__37860\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__37860\,
            I => \N__37857\
        );

    \I__9037\ : Span4Mux_v
    port map (
            O => \N__37857\,
            I => \N__37854\
        );

    \I__9036\ : Sp12to4
    port map (
            O => \N__37854\,
            I => \N__37851\
        );

    \I__9035\ : Span12Mux_h
    port map (
            O => \N__37851\,
            I => \N__37848\
        );

    \I__9034\ : Odrv12
    port map (
            O => \N__37848\,
            I => \SSEL_c\
        );

    \I__9033\ : CascadeMux
    port map (
            O => \N__37845\,
            I => \un1_bit_count_1_c1_cascade_\
        );

    \I__9032\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37839\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__37839\,
            I => \N__37836\
        );

    \I__9030\ : Span4Mux_h
    port map (
            O => \N__37836\,
            I => \N__37833\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__37833\,
            I => \OutReg_ess_RNO_1Z0Z_15\
        );

    \I__9028\ : InMux
    port map (
            O => \N__37830\,
            I => \N__37827\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__37827\,
            I => \N__37824\
        );

    \I__9026\ : Odrv12
    port map (
            O => \N__37824\,
            I => \OutReg_ess_RNO_2Z0Z_15\
        );

    \I__9025\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37818\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__37818\,
            I => \N__37815\
        );

    \I__9023\ : Odrv12
    port map (
            O => \N__37815\,
            I => \OutReg_ess_RNO_0Z0Z_15\
        );

    \I__9022\ : InMux
    port map (
            O => \N__37812\,
            I => \N__37807\
        );

    \I__9021\ : InMux
    port map (
            O => \N__37811\,
            I => \N__37802\
        );

    \I__9020\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37802\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__37807\,
            I => \N__37799\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__37802\,
            I => \bit_countZ0Z_0\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__37799\,
            I => \bit_countZ0Z_0\
        );

    \I__9016\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37791\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__37791\,
            I => \N__37788\
        );

    \I__9014\ : Span4Mux_v
    port map (
            O => \N__37788\,
            I => \N__37784\
        );

    \I__9013\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37780\
        );

    \I__9012\ : Span4Mux_h
    port map (
            O => \N__37784\,
            I => \N__37777\
        );

    \I__9011\ : InMux
    port map (
            O => \N__37783\,
            I => \N__37774\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__37780\,
            I => \N__37767\
        );

    \I__9009\ : Span4Mux_h
    port map (
            O => \N__37777\,
            I => \N__37767\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__37774\,
            I => \N__37767\
        );

    \I__9007\ : Odrv4
    port map (
            O => \N__37767\,
            I => \dataRead6_8\
        );

    \I__9006\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37756\
        );

    \I__9005\ : InMux
    port map (
            O => \N__37763\,
            I => \N__37749\
        );

    \I__9004\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37749\
        );

    \I__9003\ : InMux
    port map (
            O => \N__37761\,
            I => \N__37749\
        );

    \I__9002\ : InMux
    port map (
            O => \N__37760\,
            I => \N__37745\
        );

    \I__9001\ : InMux
    port map (
            O => \N__37759\,
            I => \N__37738\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__37756\,
            I => \N__37734\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__37749\,
            I => \N__37731\
        );

    \I__8998\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37728\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__37745\,
            I => \N__37725\
        );

    \I__8996\ : InMux
    port map (
            O => \N__37744\,
            I => \N__37722\
        );

    \I__8995\ : InMux
    port map (
            O => \N__37743\,
            I => \N__37719\
        );

    \I__8994\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37716\
        );

    \I__8993\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37713\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__37738\,
            I => \N__37709\
        );

    \I__8991\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37705\
        );

    \I__8990\ : Span4Mux_v
    port map (
            O => \N__37734\,
            I => \N__37694\
        );

    \I__8989\ : Span4Mux_h
    port map (
            O => \N__37731\,
            I => \N__37694\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__37728\,
            I => \N__37694\
        );

    \I__8987\ : Span4Mux_h
    port map (
            O => \N__37725\,
            I => \N__37689\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__37722\,
            I => \N__37689\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__37719\,
            I => \N__37686\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__37716\,
            I => \N__37681\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__37713\,
            I => \N__37681\
        );

    \I__8982\ : InMux
    port map (
            O => \N__37712\,
            I => \N__37678\
        );

    \I__8981\ : Span4Mux_h
    port map (
            O => \N__37709\,
            I => \N__37675\
        );

    \I__8980\ : InMux
    port map (
            O => \N__37708\,
            I => \N__37672\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__37705\,
            I => \N__37669\
        );

    \I__8978\ : InMux
    port map (
            O => \N__37704\,
            I => \N__37666\
        );

    \I__8977\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37663\
        );

    \I__8976\ : InMux
    port map (
            O => \N__37702\,
            I => \N__37660\
        );

    \I__8975\ : InMux
    port map (
            O => \N__37701\,
            I => \N__37657\
        );

    \I__8974\ : Span4Mux_h
    port map (
            O => \N__37694\,
            I => \N__37654\
        );

    \I__8973\ : Span4Mux_h
    port map (
            O => \N__37689\,
            I => \N__37647\
        );

    \I__8972\ : Span4Mux_h
    port map (
            O => \N__37686\,
            I => \N__37647\
        );

    \I__8971\ : Span4Mux_h
    port map (
            O => \N__37681\,
            I => \N__37647\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__37678\,
            I => \N__37640\
        );

    \I__8969\ : Span4Mux_h
    port map (
            O => \N__37675\,
            I => \N__37640\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__37672\,
            I => \N__37640\
        );

    \I__8967\ : Span12Mux_s7_v
    port map (
            O => \N__37669\,
            I => \N__37637\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__37666\,
            I => \N__37634\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__37663\,
            I => \data_receivedZ0Z_2\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__37660\,
            I => \data_receivedZ0Z_2\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__37657\,
            I => \data_receivedZ0Z_2\
        );

    \I__8962\ : Odrv4
    port map (
            O => \N__37654\,
            I => \data_receivedZ0Z_2\
        );

    \I__8961\ : Odrv4
    port map (
            O => \N__37647\,
            I => \data_receivedZ0Z_2\
        );

    \I__8960\ : Odrv4
    port map (
            O => \N__37640\,
            I => \data_receivedZ0Z_2\
        );

    \I__8959\ : Odrv12
    port map (
            O => \N__37637\,
            I => \data_receivedZ0Z_2\
        );

    \I__8958\ : Odrv4
    port map (
            O => \N__37634\,
            I => \data_receivedZ0Z_2\
        );

    \I__8957\ : CascadeMux
    port map (
            O => \N__37617\,
            I => \N__37614\
        );

    \I__8956\ : InMux
    port map (
            O => \N__37614\,
            I => \N__37609\
        );

    \I__8955\ : InMux
    port map (
            O => \N__37613\,
            I => \N__37606\
        );

    \I__8954\ : InMux
    port map (
            O => \N__37612\,
            I => \N__37603\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__37609\,
            I => \N__37600\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__37606\,
            I => \N__37595\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__37603\,
            I => \N__37595\
        );

    \I__8950\ : Span4Mux_v
    port map (
            O => \N__37600\,
            I => \N__37592\
        );

    \I__8949\ : Span4Mux_v
    port map (
            O => \N__37595\,
            I => \N__37589\
        );

    \I__8948\ : Span4Mux_h
    port map (
            O => \N__37592\,
            I => \N__37586\
        );

    \I__8947\ : Span4Mux_h
    port map (
            O => \N__37589\,
            I => \N__37583\
        );

    \I__8946\ : Odrv4
    port map (
            O => \N__37586\,
            I => \dataRead7_8\
        );

    \I__8945\ : Odrv4
    port map (
            O => \N__37583\,
            I => \dataRead7_8\
        );

    \I__8944\ : InMux
    port map (
            O => \N__37578\,
            I => \N__37575\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__37575\,
            I => \N__37572\
        );

    \I__8942\ : Odrv4
    port map (
            O => \N__37572\,
            I => \OutReg_0_4_i_m3_ns_1_8\
        );

    \I__8941\ : InMux
    port map (
            O => \N__37569\,
            I => \N__37566\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__37566\,
            I => \N__37553\
        );

    \I__8939\ : InMux
    port map (
            O => \N__37565\,
            I => \N__37550\
        );

    \I__8938\ : InMux
    port map (
            O => \N__37564\,
            I => \N__37547\
        );

    \I__8937\ : InMux
    port map (
            O => \N__37563\,
            I => \N__37544\
        );

    \I__8936\ : InMux
    port map (
            O => \N__37562\,
            I => \N__37541\
        );

    \I__8935\ : InMux
    port map (
            O => \N__37561\,
            I => \N__37538\
        );

    \I__8934\ : InMux
    port map (
            O => \N__37560\,
            I => \N__37534\
        );

    \I__8933\ : InMux
    port map (
            O => \N__37559\,
            I => \N__37531\
        );

    \I__8932\ : InMux
    port map (
            O => \N__37558\,
            I => \N__37528\
        );

    \I__8931\ : InMux
    port map (
            O => \N__37557\,
            I => \N__37525\
        );

    \I__8930\ : InMux
    port map (
            O => \N__37556\,
            I => \N__37522\
        );

    \I__8929\ : Span4Mux_h
    port map (
            O => \N__37553\,
            I => \N__37514\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__37550\,
            I => \N__37514\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__37547\,
            I => \N__37514\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__37544\,
            I => \N__37508\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__37541\,
            I => \N__37499\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__37538\,
            I => \N__37496\
        );

    \I__8923\ : InMux
    port map (
            O => \N__37537\,
            I => \N__37493\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__37534\,
            I => \N__37486\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__37531\,
            I => \N__37486\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__37528\,
            I => \N__37486\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__37525\,
            I => \N__37483\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__37522\,
            I => \N__37480\
        );

    \I__8917\ : InMux
    port map (
            O => \N__37521\,
            I => \N__37477\
        );

    \I__8916\ : Span4Mux_v
    port map (
            O => \N__37514\,
            I => \N__37474\
        );

    \I__8915\ : InMux
    port map (
            O => \N__37513\,
            I => \N__37469\
        );

    \I__8914\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37469\
        );

    \I__8913\ : InMux
    port map (
            O => \N__37511\,
            I => \N__37466\
        );

    \I__8912\ : Span12Mux_v
    port map (
            O => \N__37508\,
            I => \N__37463\
        );

    \I__8911\ : InMux
    port map (
            O => \N__37507\,
            I => \N__37456\
        );

    \I__8910\ : InMux
    port map (
            O => \N__37506\,
            I => \N__37456\
        );

    \I__8909\ : InMux
    port map (
            O => \N__37505\,
            I => \N__37456\
        );

    \I__8908\ : InMux
    port map (
            O => \N__37504\,
            I => \N__37449\
        );

    \I__8907\ : InMux
    port map (
            O => \N__37503\,
            I => \N__37449\
        );

    \I__8906\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37449\
        );

    \I__8905\ : Span4Mux_h
    port map (
            O => \N__37499\,
            I => \N__37444\
        );

    \I__8904\ : Span4Mux_h
    port map (
            O => \N__37496\,
            I => \N__37444\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__37493\,
            I => \N__37439\
        );

    \I__8902\ : Span4Mux_h
    port map (
            O => \N__37486\,
            I => \N__37439\
        );

    \I__8901\ : Span4Mux_h
    port map (
            O => \N__37483\,
            I => \N__37434\
        );

    \I__8900\ : Span4Mux_h
    port map (
            O => \N__37480\,
            I => \N__37434\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__37477\,
            I => \N__37427\
        );

    \I__8898\ : Span4Mux_h
    port map (
            O => \N__37474\,
            I => \N__37427\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__37469\,
            I => \N__37427\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__37466\,
            I => \data_receivedZ0Z_1\
        );

    \I__8895\ : Odrv12
    port map (
            O => \N__37463\,
            I => \data_receivedZ0Z_1\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__37456\,
            I => \data_receivedZ0Z_1\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__37449\,
            I => \data_receivedZ0Z_1\
        );

    \I__8892\ : Odrv4
    port map (
            O => \N__37444\,
            I => \data_receivedZ0Z_1\
        );

    \I__8891\ : Odrv4
    port map (
            O => \N__37439\,
            I => \data_receivedZ0Z_1\
        );

    \I__8890\ : Odrv4
    port map (
            O => \N__37434\,
            I => \data_receivedZ0Z_1\
        );

    \I__8889\ : Odrv4
    port map (
            O => \N__37427\,
            I => \data_receivedZ0Z_1\
        );

    \I__8888\ : CascadeMux
    port map (
            O => \N__37410\,
            I => \OutReg_esr_RNO_1Z0Z_8_cascade_\
        );

    \I__8887\ : InMux
    port map (
            O => \N__37407\,
            I => \N__37404\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__37404\,
            I => \N__37401\
        );

    \I__8885\ : Odrv12
    port map (
            O => \N__37401\,
            I => \OutRegZ0Z_7\
        );

    \I__8884\ : CascadeMux
    port map (
            O => \N__37398\,
            I => \OutReg_esr_RNO_0Z0Z_8_cascade_\
        );

    \I__8883\ : InMux
    port map (
            O => \N__37395\,
            I => \N__37389\
        );

    \I__8882\ : InMux
    port map (
            O => \N__37394\,
            I => \N__37389\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__37389\,
            I => \N__37382\
        );

    \I__8880\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37375\
        );

    \I__8879\ : InMux
    port map (
            O => \N__37387\,
            I => \N__37371\
        );

    \I__8878\ : InMux
    port map (
            O => \N__37386\,
            I => \N__37366\
        );

    \I__8877\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37366\
        );

    \I__8876\ : Span4Mux_h
    port map (
            O => \N__37382\,
            I => \N__37363\
        );

    \I__8875\ : InMux
    port map (
            O => \N__37381\,
            I => \N__37360\
        );

    \I__8874\ : InMux
    port map (
            O => \N__37380\,
            I => \N__37357\
        );

    \I__8873\ : InMux
    port map (
            O => \N__37379\,
            I => \N__37352\
        );

    \I__8872\ : InMux
    port map (
            O => \N__37378\,
            I => \N__37352\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__37375\,
            I => \N__37348\
        );

    \I__8870\ : InMux
    port map (
            O => \N__37374\,
            I => \N__37345\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__37371\,
            I => \N__37341\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__37366\,
            I => \N__37338\
        );

    \I__8867\ : Span4Mux_h
    port map (
            O => \N__37363\,
            I => \N__37333\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__37360\,
            I => \N__37333\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__37357\,
            I => \N__37327\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__37352\,
            I => \N__37327\
        );

    \I__8863\ : InMux
    port map (
            O => \N__37351\,
            I => \N__37324\
        );

    \I__8862\ : Span4Mux_v
    port map (
            O => \N__37348\,
            I => \N__37317\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__37345\,
            I => \N__37317\
        );

    \I__8860\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37314\
        );

    \I__8859\ : Span4Mux_h
    port map (
            O => \N__37341\,
            I => \N__37307\
        );

    \I__8858\ : Span4Mux_h
    port map (
            O => \N__37338\,
            I => \N__37307\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__37333\,
            I => \N__37304\
        );

    \I__8856\ : InMux
    port map (
            O => \N__37332\,
            I => \N__37301\
        );

    \I__8855\ : Span4Mux_v
    port map (
            O => \N__37327\,
            I => \N__37296\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__37324\,
            I => \N__37296\
        );

    \I__8853\ : InMux
    port map (
            O => \N__37323\,
            I => \N__37293\
        );

    \I__8852\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37290\
        );

    \I__8851\ : Span4Mux_h
    port map (
            O => \N__37317\,
            I => \N__37285\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__37314\,
            I => \N__37285\
        );

    \I__8849\ : InMux
    port map (
            O => \N__37313\,
            I => \N__37280\
        );

    \I__8848\ : InMux
    port map (
            O => \N__37312\,
            I => \N__37280\
        );

    \I__8847\ : Odrv4
    port map (
            O => \N__37307\,
            I => \un1_OutReg51_4_0_i_o3_2\
        );

    \I__8846\ : Odrv4
    port map (
            O => \N__37304\,
            I => \un1_OutReg51_4_0_i_o3_2\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__37301\,
            I => \un1_OutReg51_4_0_i_o3_2\
        );

    \I__8844\ : Odrv4
    port map (
            O => \N__37296\,
            I => \un1_OutReg51_4_0_i_o3_2\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__37293\,
            I => \un1_OutReg51_4_0_i_o3_2\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__37290\,
            I => \un1_OutReg51_4_0_i_o3_2\
        );

    \I__8841\ : Odrv4
    port map (
            O => \N__37285\,
            I => \un1_OutReg51_4_0_i_o3_2\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__37280\,
            I => \un1_OutReg51_4_0_i_o3_2\
        );

    \I__8839\ : InMux
    port map (
            O => \N__37263\,
            I => \N__37260\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__37260\,
            I => \N__37257\
        );

    \I__8837\ : Sp12to4
    port map (
            O => \N__37257\,
            I => \N__37254\
        );

    \I__8836\ : Odrv12
    port map (
            O => \N__37254\,
            I => \OutRegZ0Z_8\
        );

    \I__8835\ : CEMux
    port map (
            O => \N__37251\,
            I => \N__37247\
        );

    \I__8834\ : CEMux
    port map (
            O => \N__37250\,
            I => \N__37237\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__37247\,
            I => \N__37234\
        );

    \I__8832\ : CEMux
    port map (
            O => \N__37246\,
            I => \N__37231\
        );

    \I__8831\ : CEMux
    port map (
            O => \N__37245\,
            I => \N__37228\
        );

    \I__8830\ : CEMux
    port map (
            O => \N__37244\,
            I => \N__37225\
        );

    \I__8829\ : CEMux
    port map (
            O => \N__37243\,
            I => \N__37221\
        );

    \I__8828\ : CEMux
    port map (
            O => \N__37242\,
            I => \N__37218\
        );

    \I__8827\ : CEMux
    port map (
            O => \N__37241\,
            I => \N__37215\
        );

    \I__8826\ : CEMux
    port map (
            O => \N__37240\,
            I => \N__37212\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__37237\,
            I => \N__37207\
        );

    \I__8824\ : Span4Mux_h
    port map (
            O => \N__37234\,
            I => \N__37202\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__37231\,
            I => \N__37202\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__37228\,
            I => \N__37197\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__37225\,
            I => \N__37197\
        );

    \I__8820\ : CEMux
    port map (
            O => \N__37224\,
            I => \N__37194\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__37221\,
            I => \N__37191\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__37218\,
            I => \N__37186\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__37215\,
            I => \N__37186\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__37212\,
            I => \N__37183\
        );

    \I__8815\ : CEMux
    port map (
            O => \N__37211\,
            I => \N__37180\
        );

    \I__8814\ : CEMux
    port map (
            O => \N__37210\,
            I => \N__37177\
        );

    \I__8813\ : Span4Mux_h
    port map (
            O => \N__37207\,
            I => \N__37174\
        );

    \I__8812\ : Span4Mux_v
    port map (
            O => \N__37202\,
            I => \N__37171\
        );

    \I__8811\ : Span4Mux_h
    port map (
            O => \N__37197\,
            I => \N__37168\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__37194\,
            I => \N__37165\
        );

    \I__8809\ : Span4Mux_v
    port map (
            O => \N__37191\,
            I => \N__37160\
        );

    \I__8808\ : Span4Mux_h
    port map (
            O => \N__37186\,
            I => \N__37160\
        );

    \I__8807\ : Sp12to4
    port map (
            O => \N__37183\,
            I => \N__37155\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__37180\,
            I => \N__37155\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__37177\,
            I => \N__37152\
        );

    \I__8804\ : Odrv4
    port map (
            O => \N__37174\,
            I => \N_863_0\
        );

    \I__8803\ : Odrv4
    port map (
            O => \N__37171\,
            I => \N_863_0\
        );

    \I__8802\ : Odrv4
    port map (
            O => \N__37168\,
            I => \N_863_0\
        );

    \I__8801\ : Odrv4
    port map (
            O => \N__37165\,
            I => \N_863_0\
        );

    \I__8800\ : Odrv4
    port map (
            O => \N__37160\,
            I => \N_863_0\
        );

    \I__8799\ : Odrv12
    port map (
            O => \N__37155\,
            I => \N_863_0\
        );

    \I__8798\ : Odrv12
    port map (
            O => \N__37152\,
            I => \N_863_0\
        );

    \I__8797\ : SRMux
    port map (
            O => \N__37137\,
            I => \N__37125\
        );

    \I__8796\ : SRMux
    port map (
            O => \N__37136\,
            I => \N__37122\
        );

    \I__8795\ : SRMux
    port map (
            O => \N__37135\,
            I => \N__37119\
        );

    \I__8794\ : SRMux
    port map (
            O => \N__37134\,
            I => \N__37116\
        );

    \I__8793\ : SRMux
    port map (
            O => \N__37133\,
            I => \N__37112\
        );

    \I__8792\ : SRMux
    port map (
            O => \N__37132\,
            I => \N__37109\
        );

    \I__8791\ : SRMux
    port map (
            O => \N__37131\,
            I => \N__37106\
        );

    \I__8790\ : SRMux
    port map (
            O => \N__37130\,
            I => \N__37103\
        );

    \I__8789\ : SRMux
    port map (
            O => \N__37129\,
            I => \N__37100\
        );

    \I__8788\ : SRMux
    port map (
            O => \N__37128\,
            I => \N__37096\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__37125\,
            I => \N__37093\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__37122\,
            I => \N__37090\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__37119\,
            I => \N__37087\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__37116\,
            I => \N__37084\
        );

    \I__8783\ : SRMux
    port map (
            O => \N__37115\,
            I => \N__37081\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__37112\,
            I => \N__37078\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__37109\,
            I => \N__37075\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__37106\,
            I => \N__37072\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__37103\,
            I => \N__37067\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__37100\,
            I => \N__37067\
        );

    \I__8777\ : SRMux
    port map (
            O => \N__37099\,
            I => \N__37064\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__37096\,
            I => \N__37061\
        );

    \I__8775\ : Span4Mux_h
    port map (
            O => \N__37093\,
            I => \N__37055\
        );

    \I__8774\ : Span4Mux_h
    port map (
            O => \N__37090\,
            I => \N__37055\
        );

    \I__8773\ : Span4Mux_v
    port map (
            O => \N__37087\,
            I => \N__37050\
        );

    \I__8772\ : Span4Mux_h
    port map (
            O => \N__37084\,
            I => \N__37050\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__37081\,
            I => \N__37047\
        );

    \I__8770\ : Span4Mux_h
    port map (
            O => \N__37078\,
            I => \N__37038\
        );

    \I__8769\ : Span4Mux_v
    port map (
            O => \N__37075\,
            I => \N__37038\
        );

    \I__8768\ : Span4Mux_v
    port map (
            O => \N__37072\,
            I => \N__37038\
        );

    \I__8767\ : Span4Mux_h
    port map (
            O => \N__37067\,
            I => \N__37038\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__37064\,
            I => \N__37033\
        );

    \I__8765\ : Span4Mux_h
    port map (
            O => \N__37061\,
            I => \N__37033\
        );

    \I__8764\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37030\
        );

    \I__8763\ : Odrv4
    port map (
            O => \N__37055\,
            I => \OutReg_0_sqmuxa\
        );

    \I__8762\ : Odrv4
    port map (
            O => \N__37050\,
            I => \OutReg_0_sqmuxa\
        );

    \I__8761\ : Odrv4
    port map (
            O => \N__37047\,
            I => \OutReg_0_sqmuxa\
        );

    \I__8760\ : Odrv4
    port map (
            O => \N__37038\,
            I => \OutReg_0_sqmuxa\
        );

    \I__8759\ : Odrv4
    port map (
            O => \N__37033\,
            I => \OutReg_0_sqmuxa\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__37030\,
            I => \OutReg_0_sqmuxa\
        );

    \I__8757\ : InMux
    port map (
            O => \N__37017\,
            I => \N__37014\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__37014\,
            I => \N__37009\
        );

    \I__8755\ : InMux
    port map (
            O => \N__37013\,
            I => \N__37006\
        );

    \I__8754\ : InMux
    port map (
            O => \N__37012\,
            I => \N__37003\
        );

    \I__8753\ : Span4Mux_v
    port map (
            O => \N__37009\,
            I => \N__37000\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__37006\,
            I => \N__36995\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__37003\,
            I => \N__36995\
        );

    \I__8750\ : Sp12to4
    port map (
            O => \N__37000\,
            I => \N__36992\
        );

    \I__8749\ : Span4Mux_h
    port map (
            O => \N__36995\,
            I => \N__36989\
        );

    \I__8748\ : Odrv12
    port map (
            O => \N__36992\,
            I => \dataRead1_8\
        );

    \I__8747\ : Odrv4
    port map (
            O => \N__36989\,
            I => \dataRead1_8\
        );

    \I__8746\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36981\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__36981\,
            I => \N__36977\
        );

    \I__8744\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36974\
        );

    \I__8743\ : Span4Mux_v
    port map (
            O => \N__36977\,
            I => \N__36970\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__36974\,
            I => \N__36967\
        );

    \I__8741\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36964\
        );

    \I__8740\ : Span4Mux_h
    port map (
            O => \N__36970\,
            I => \N__36961\
        );

    \I__8739\ : Span12Mux_h
    port map (
            O => \N__36967\,
            I => \N__36958\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__36964\,
            I => \N__36955\
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__36961\,
            I => \dataRead5_8\
        );

    \I__8736\ : Odrv12
    port map (
            O => \N__36958\,
            I => \dataRead5_8\
        );

    \I__8735\ : Odrv4
    port map (
            O => \N__36955\,
            I => \dataRead5_8\
        );

    \I__8734\ : IoInMux
    port map (
            O => \N__36948\,
            I => \N__36945\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__36945\,
            I => \PWM3_obufLegalizeSB_DFFNet\
        );

    \I__8732\ : IoInMux
    port map (
            O => \N__36942\,
            I => \N__36939\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__36939\,
            I => \MISO_obufLegalizeSB_DFFNet\
        );

    \I__8730\ : ClkMux
    port map (
            O => \N__36936\,
            I => \N__36933\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__36933\,
            I => \N__36929\
        );

    \I__8728\ : ClkMux
    port map (
            O => \N__36932\,
            I => \N__36926\
        );

    \I__8727\ : Span4Mux_h
    port map (
            O => \N__36929\,
            I => \N__36920\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__36926\,
            I => \N__36920\
        );

    \I__8725\ : ClkMux
    port map (
            O => \N__36925\,
            I => \N__36917\
        );

    \I__8724\ : Span4Mux_h
    port map (
            O => \N__36920\,
            I => \N__36913\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__36917\,
            I => \N__36910\
        );

    \I__8722\ : ClkMux
    port map (
            O => \N__36916\,
            I => \N__36907\
        );

    \I__8721\ : Span4Mux_h
    port map (
            O => \N__36913\,
            I => \N__36899\
        );

    \I__8720\ : Span4Mux_h
    port map (
            O => \N__36910\,
            I => \N__36899\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__36907\,
            I => \N__36899\
        );

    \I__8718\ : ClkMux
    port map (
            O => \N__36906\,
            I => \N__36896\
        );

    \I__8717\ : Sp12to4
    port map (
            O => \N__36899\,
            I => \N__36893\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__36896\,
            I => \N__36890\
        );

    \I__8715\ : Span12Mux_h
    port map (
            O => \N__36893\,
            I => \N__36887\
        );

    \I__8714\ : Span4Mux_h
    port map (
            O => \N__36890\,
            I => \N__36884\
        );

    \I__8713\ : Span12Mux_v
    port map (
            O => \N__36887\,
            I => \N__36881\
        );

    \I__8712\ : Span4Mux_h
    port map (
            O => \N__36884\,
            I => \N__36878\
        );

    \I__8711\ : Odrv12
    port map (
            O => \N__36881\,
            I => \internalOscilatorOutputNet\
        );

    \I__8710\ : Odrv4
    port map (
            O => \N__36878\,
            I => \internalOscilatorOutputNet\
        );

    \I__8709\ : InMux
    port map (
            O => \N__36873\,
            I => \N__36868\
        );

    \I__8708\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36865\
        );

    \I__8707\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36862\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36859\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__36865\,
            I => \N__36856\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36853\
        );

    \I__8703\ : Span4Mux_v
    port map (
            O => \N__36859\,
            I => \N__36850\
        );

    \I__8702\ : Span4Mux_h
    port map (
            O => \N__36856\,
            I => \N__36847\
        );

    \I__8701\ : Span4Mux_h
    port map (
            O => \N__36853\,
            I => \N__36844\
        );

    \I__8700\ : Span4Mux_h
    port map (
            O => \N__36850\,
            I => \N__36841\
        );

    \I__8699\ : Sp12to4
    port map (
            O => \N__36847\,
            I => \N__36838\
        );

    \I__8698\ : Odrv4
    port map (
            O => \N__36844\,
            I => \dataRead5_5\
        );

    \I__8697\ : Odrv4
    port map (
            O => \N__36841\,
            I => \dataRead5_5\
        );

    \I__8696\ : Odrv12
    port map (
            O => \N__36838\,
            I => \dataRead5_5\
        );

    \I__8695\ : CascadeMux
    port map (
            O => \N__36831\,
            I => \N__36828\
        );

    \I__8694\ : InMux
    port map (
            O => \N__36828\,
            I => \N__36824\
        );

    \I__8693\ : InMux
    port map (
            O => \N__36827\,
            I => \N__36821\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__36824\,
            I => \N__36818\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__36821\,
            I => \N__36814\
        );

    \I__8690\ : Span4Mux_h
    port map (
            O => \N__36818\,
            I => \N__36811\
        );

    \I__8689\ : InMux
    port map (
            O => \N__36817\,
            I => \N__36808\
        );

    \I__8688\ : Span4Mux_v
    port map (
            O => \N__36814\,
            I => \N__36805\
        );

    \I__8687\ : Span4Mux_h
    port map (
            O => \N__36811\,
            I => \N__36800\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__36808\,
            I => \N__36800\
        );

    \I__8685\ : Odrv4
    port map (
            O => \N__36805\,
            I => \dataRead1_5\
        );

    \I__8684\ : Odrv4
    port map (
            O => \N__36800\,
            I => \dataRead1_5\
        );

    \I__8683\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36792\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__36792\,
            I => \N__36789\
        );

    \I__8681\ : Span4Mux_v
    port map (
            O => \N__36789\,
            I => \N__36786\
        );

    \I__8680\ : Odrv4
    port map (
            O => \N__36786\,
            I => \OutReg_0_5_i_m3_ns_1_5\
        );

    \I__8679\ : InMux
    port map (
            O => \N__36783\,
            I => \N__36780\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__36780\,
            I => \N__36777\
        );

    \I__8677\ : Span4Mux_v
    port map (
            O => \N__36777\,
            I => \N__36773\
        );

    \I__8676\ : InMux
    port map (
            O => \N__36776\,
            I => \N__36770\
        );

    \I__8675\ : Span4Mux_h
    port map (
            O => \N__36773\,
            I => \N__36767\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__36770\,
            I => \N__36763\
        );

    \I__8673\ : Span4Mux_h
    port map (
            O => \N__36767\,
            I => \N__36760\
        );

    \I__8672\ : InMux
    port map (
            O => \N__36766\,
            I => \N__36757\
        );

    \I__8671\ : Odrv12
    port map (
            O => \N__36763\,
            I => \dataRead6_5\
        );

    \I__8670\ : Odrv4
    port map (
            O => \N__36760\,
            I => \dataRead6_5\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__36757\,
            I => \dataRead6_5\
        );

    \I__8668\ : CascadeMux
    port map (
            O => \N__36750\,
            I => \N__36747\
        );

    \I__8667\ : InMux
    port map (
            O => \N__36747\,
            I => \N__36743\
        );

    \I__8666\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36740\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__36743\,
            I => \N__36736\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__36740\,
            I => \N__36733\
        );

    \I__8663\ : InMux
    port map (
            O => \N__36739\,
            I => \N__36730\
        );

    \I__8662\ : Span4Mux_v
    port map (
            O => \N__36736\,
            I => \N__36727\
        );

    \I__8661\ : Span4Mux_h
    port map (
            O => \N__36733\,
            I => \N__36722\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__36730\,
            I => \N__36722\
        );

    \I__8659\ : Span4Mux_h
    port map (
            O => \N__36727\,
            I => \N__36719\
        );

    \I__8658\ : Span4Mux_v
    port map (
            O => \N__36722\,
            I => \N__36716\
        );

    \I__8657\ : Odrv4
    port map (
            O => \N__36719\,
            I => \dataRead7_5\
        );

    \I__8656\ : Odrv4
    port map (
            O => \N__36716\,
            I => \dataRead7_5\
        );

    \I__8655\ : InMux
    port map (
            O => \N__36711\,
            I => \N__36708\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__36708\,
            I => \N__36705\
        );

    \I__8653\ : Span4Mux_v
    port map (
            O => \N__36705\,
            I => \N__36702\
        );

    \I__8652\ : Span4Mux_h
    port map (
            O => \N__36702\,
            I => \N__36699\
        );

    \I__8651\ : Odrv4
    port map (
            O => \N__36699\,
            I => \OutReg_0_4_i_m3_ns_1_5\
        );

    \I__8650\ : CascadeMux
    port map (
            O => \N__36696\,
            I => \OutReg_ess_RNO_1Z0Z_5_cascade_\
        );

    \I__8649\ : InMux
    port map (
            O => \N__36693\,
            I => \N__36690\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__36690\,
            I => \OutReg_ess_RNO_2Z0Z_5\
        );

    \I__8647\ : InMux
    port map (
            O => \N__36687\,
            I => \N__36684\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__36684\,
            I => \OutReg_ess_RNO_0Z0Z_5\
        );

    \I__8645\ : CascadeMux
    port map (
            O => \N__36681\,
            I => \N__36678\
        );

    \I__8644\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36675\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__36675\,
            I => \N__36672\
        );

    \I__8642\ : Span4Mux_h
    port map (
            O => \N__36672\,
            I => \N__36669\
        );

    \I__8641\ : Odrv4
    port map (
            O => \N__36669\,
            I => \OutRegZ0Z_4\
        );

    \I__8640\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36663\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__36663\,
            I => \N__36660\
        );

    \I__8638\ : Span4Mux_h
    port map (
            O => \N__36660\,
            I => \N__36657\
        );

    \I__8637\ : Odrv4
    port map (
            O => \N__36657\,
            I => \OutRegZ0Z_5\
        );

    \I__8636\ : InMux
    port map (
            O => \N__36654\,
            I => \N__36651\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__36651\,
            I => \N__36648\
        );

    \I__8634\ : Span4Mux_h
    port map (
            O => \N__36648\,
            I => \N__36645\
        );

    \I__8633\ : Odrv4
    port map (
            O => \N__36645\,
            I => \OutRegZ0Z_15\
        );

    \I__8632\ : CascadeMux
    port map (
            O => \N__36642\,
            I => \dataOut_RNOZ0Z_0_cascade_\
        );

    \I__8631\ : IoInMux
    port map (
            O => \N__36639\,
            I => \N__36636\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__36636\,
            I => \N__36633\
        );

    \I__8629\ : Span4Mux_s2_v
    port map (
            O => \N__36633\,
            I => \N__36630\
        );

    \I__8628\ : Span4Mux_v
    port map (
            O => \N__36630\,
            I => \N__36626\
        );

    \I__8627\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36623\
        );

    \I__8626\ : Odrv4
    port map (
            O => \N__36626\,
            I => \MISO_c\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__36623\,
            I => \MISO_c\
        );

    \I__8624\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36613\
        );

    \I__8623\ : InMux
    port map (
            O => \N__36617\,
            I => \N__36610\
        );

    \I__8622\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36607\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__36613\,
            I => \N__36604\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__36610\,
            I => \PWMInstance2.periodCounterZ0Z_14\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__36607\,
            I => \PWMInstance2.periodCounterZ0Z_14\
        );

    \I__8618\ : Odrv4
    port map (
            O => \N__36604\,
            I => \PWMInstance2.periodCounterZ0Z_14\
        );

    \I__8617\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36592\
        );

    \I__8616\ : InMux
    port map (
            O => \N__36596\,
            I => \N__36589\
        );

    \I__8615\ : InMux
    port map (
            O => \N__36595\,
            I => \N__36586\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__36592\,
            I => \N__36581\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__36589\,
            I => \N__36581\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__36586\,
            I => \PWMInstance2.periodCounterZ0Z_2\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__36581\,
            I => \PWMInstance2.periodCounterZ0Z_2\
        );

    \I__8610\ : InMux
    port map (
            O => \N__36576\,
            I => \N__36569\
        );

    \I__8609\ : InMux
    port map (
            O => \N__36575\,
            I => \N__36569\
        );

    \I__8608\ : InMux
    port map (
            O => \N__36574\,
            I => \N__36566\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__36569\,
            I => \N__36563\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__36566\,
            I => \PWMInstance2.periodCounterZ0Z_4\
        );

    \I__8605\ : Odrv4
    port map (
            O => \N__36563\,
            I => \PWMInstance2.periodCounterZ0Z_4\
        );

    \I__8604\ : InMux
    port map (
            O => \N__36558\,
            I => \N__36553\
        );

    \I__8603\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36550\
        );

    \I__8602\ : InMux
    port map (
            O => \N__36556\,
            I => \N__36547\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__36553\,
            I => \N__36544\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__36550\,
            I => \PWMInstance2.periodCounterZ0Z_12\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__36547\,
            I => \PWMInstance2.periodCounterZ0Z_12\
        );

    \I__8598\ : Odrv4
    port map (
            O => \N__36544\,
            I => \PWMInstance2.periodCounterZ0Z_12\
        );

    \I__8597\ : CascadeMux
    port map (
            O => \N__36537\,
            I => \PWMInstance2.un1_periodCounter12_1_0_a2_0_0_cascade_\
        );

    \I__8596\ : InMux
    port map (
            O => \N__36534\,
            I => \N__36531\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__36531\,
            I => \N__36528\
        );

    \I__8594\ : Odrv4
    port map (
            O => \N__36528\,
            I => \PWMInstance2.un1_periodCounter12_1_0_a2_0_12\
        );

    \I__8593\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36522\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__36522\,
            I => \N__36518\
        );

    \I__8591\ : InMux
    port map (
            O => \N__36521\,
            I => \N__36515\
        );

    \I__8590\ : Span4Mux_s2_v
    port map (
            O => \N__36518\,
            I => \N__36507\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__36515\,
            I => \N__36507\
        );

    \I__8588\ : InMux
    port map (
            O => \N__36514\,
            I => \N__36504\
        );

    \I__8587\ : InMux
    port map (
            O => \N__36513\,
            I => \N__36498\
        );

    \I__8586\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36495\
        );

    \I__8585\ : Span4Mux_h
    port map (
            O => \N__36507\,
            I => \N__36489\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__36504\,
            I => \N__36489\
        );

    \I__8583\ : InMux
    port map (
            O => \N__36503\,
            I => \N__36480\
        );

    \I__8582\ : InMux
    port map (
            O => \N__36502\,
            I => \N__36477\
        );

    \I__8581\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36474\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__36498\,
            I => \N__36471\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__36495\,
            I => \N__36468\
        );

    \I__8578\ : InMux
    port map (
            O => \N__36494\,
            I => \N__36465\
        );

    \I__8577\ : Span4Mux_v
    port map (
            O => \N__36489\,
            I => \N__36462\
        );

    \I__8576\ : InMux
    port map (
            O => \N__36488\,
            I => \N__36451\
        );

    \I__8575\ : InMux
    port map (
            O => \N__36487\,
            I => \N__36451\
        );

    \I__8574\ : InMux
    port map (
            O => \N__36486\,
            I => \N__36451\
        );

    \I__8573\ : InMux
    port map (
            O => \N__36485\,
            I => \N__36451\
        );

    \I__8572\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36451\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__36483\,
            I => \N__36448\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__36480\,
            I => \N__36445\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__36477\,
            I => \N__36442\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__36474\,
            I => \N__36439\
        );

    \I__8567\ : Span4Mux_v
    port map (
            O => \N__36471\,
            I => \N__36435\
        );

    \I__8566\ : Span4Mux_v
    port map (
            O => \N__36468\,
            I => \N__36430\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__36465\,
            I => \N__36430\
        );

    \I__8564\ : Span4Mux_h
    port map (
            O => \N__36462\,
            I => \N__36427\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__36451\,
            I => \N__36424\
        );

    \I__8562\ : InMux
    port map (
            O => \N__36448\,
            I => \N__36421\
        );

    \I__8561\ : Span12Mux_h
    port map (
            O => \N__36445\,
            I => \N__36418\
        );

    \I__8560\ : Span4Mux_v
    port map (
            O => \N__36442\,
            I => \N__36415\
        );

    \I__8559\ : Span4Mux_v
    port map (
            O => \N__36439\,
            I => \N__36412\
        );

    \I__8558\ : InMux
    port map (
            O => \N__36438\,
            I => \N__36409\
        );

    \I__8557\ : Span4Mux_h
    port map (
            O => \N__36435\,
            I => \N__36402\
        );

    \I__8556\ : Span4Mux_v
    port map (
            O => \N__36430\,
            I => \N__36402\
        );

    \I__8555\ : Span4Mux_v
    port map (
            O => \N__36427\,
            I => \N__36402\
        );

    \I__8554\ : Span4Mux_v
    port map (
            O => \N__36424\,
            I => \N__36397\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__36421\,
            I => \N__36397\
        );

    \I__8552\ : Odrv12
    port map (
            O => \N__36418\,
            I => \dataWriteZ0Z_4\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__36415\,
            I => \dataWriteZ0Z_4\
        );

    \I__8550\ : Odrv4
    port map (
            O => \N__36412\,
            I => \dataWriteZ0Z_4\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__36409\,
            I => \dataWriteZ0Z_4\
        );

    \I__8548\ : Odrv4
    port map (
            O => \N__36402\,
            I => \dataWriteZ0Z_4\
        );

    \I__8547\ : Odrv4
    port map (
            O => \N__36397\,
            I => \dataWriteZ0Z_4\
        );

    \I__8546\ : InMux
    port map (
            O => \N__36384\,
            I => \N__36381\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__36381\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_4\
        );

    \I__8544\ : CascadeMux
    port map (
            O => \N__36378\,
            I => \N__36373\
        );

    \I__8543\ : InMux
    port map (
            O => \N__36377\,
            I => \N__36363\
        );

    \I__8542\ : InMux
    port map (
            O => \N__36376\,
            I => \N__36359\
        );

    \I__8541\ : InMux
    port map (
            O => \N__36373\,
            I => \N__36348\
        );

    \I__8540\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36348\
        );

    \I__8539\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36348\
        );

    \I__8538\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36348\
        );

    \I__8537\ : InMux
    port map (
            O => \N__36369\,
            I => \N__36348\
        );

    \I__8536\ : InMux
    port map (
            O => \N__36368\,
            I => \N__36342\
        );

    \I__8535\ : InMux
    port map (
            O => \N__36367\,
            I => \N__36339\
        );

    \I__8534\ : InMux
    port map (
            O => \N__36366\,
            I => \N__36336\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__36363\,
            I => \N__36333\
        );

    \I__8532\ : InMux
    port map (
            O => \N__36362\,
            I => \N__36329\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__36359\,
            I => \N__36326\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__36348\,
            I => \N__36323\
        );

    \I__8529\ : InMux
    port map (
            O => \N__36347\,
            I => \N__36320\
        );

    \I__8528\ : InMux
    port map (
            O => \N__36346\,
            I => \N__36317\
        );

    \I__8527\ : InMux
    port map (
            O => \N__36345\,
            I => \N__36314\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__36342\,
            I => \N__36311\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__36339\,
            I => \N__36308\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__36336\,
            I => \N__36305\
        );

    \I__8523\ : Span4Mux_v
    port map (
            O => \N__36333\,
            I => \N__36302\
        );

    \I__8522\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36299\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__36329\,
            I => \N__36296\
        );

    \I__8520\ : Span4Mux_v
    port map (
            O => \N__36326\,
            I => \N__36293\
        );

    \I__8519\ : Span4Mux_v
    port map (
            O => \N__36323\,
            I => \N__36290\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__36320\,
            I => \N__36285\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__36317\,
            I => \N__36285\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__36314\,
            I => \N__36281\
        );

    \I__8515\ : Span4Mux_v
    port map (
            O => \N__36311\,
            I => \N__36278\
        );

    \I__8514\ : Span4Mux_v
    port map (
            O => \N__36308\,
            I => \N__36271\
        );

    \I__8513\ : Span4Mux_v
    port map (
            O => \N__36305\,
            I => \N__36271\
        );

    \I__8512\ : Span4Mux_v
    port map (
            O => \N__36302\,
            I => \N__36271\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__36299\,
            I => \N__36266\
        );

    \I__8510\ : Span4Mux_v
    port map (
            O => \N__36296\,
            I => \N__36266\
        );

    \I__8509\ : Span4Mux_h
    port map (
            O => \N__36293\,
            I => \N__36263\
        );

    \I__8508\ : Span4Mux_h
    port map (
            O => \N__36290\,
            I => \N__36260\
        );

    \I__8507\ : Span4Mux_h
    port map (
            O => \N__36285\,
            I => \N__36257\
        );

    \I__8506\ : InMux
    port map (
            O => \N__36284\,
            I => \N__36254\
        );

    \I__8505\ : Span4Mux_h
    port map (
            O => \N__36281\,
            I => \N__36251\
        );

    \I__8504\ : Span4Mux_v
    port map (
            O => \N__36278\,
            I => \N__36246\
        );

    \I__8503\ : Span4Mux_h
    port map (
            O => \N__36271\,
            I => \N__36246\
        );

    \I__8502\ : Span4Mux_v
    port map (
            O => \N__36266\,
            I => \N__36239\
        );

    \I__8501\ : Span4Mux_h
    port map (
            O => \N__36263\,
            I => \N__36239\
        );

    \I__8500\ : Span4Mux_v
    port map (
            O => \N__36260\,
            I => \N__36239\
        );

    \I__8499\ : Span4Mux_v
    port map (
            O => \N__36257\,
            I => \N__36236\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__36254\,
            I => \dataWriteZ0Z_5\
        );

    \I__8497\ : Odrv4
    port map (
            O => \N__36251\,
            I => \dataWriteZ0Z_5\
        );

    \I__8496\ : Odrv4
    port map (
            O => \N__36246\,
            I => \dataWriteZ0Z_5\
        );

    \I__8495\ : Odrv4
    port map (
            O => \N__36239\,
            I => \dataWriteZ0Z_5\
        );

    \I__8494\ : Odrv4
    port map (
            O => \N__36236\,
            I => \dataWriteZ0Z_5\
        );

    \I__8493\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36222\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__36222\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_5\
        );

    \I__8491\ : InMux
    port map (
            O => \N__36219\,
            I => \N__36212\
        );

    \I__8490\ : InMux
    port map (
            O => \N__36218\,
            I => \N__36212\
        );

    \I__8489\ : InMux
    port map (
            O => \N__36217\,
            I => \N__36209\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__36212\,
            I => \N__36206\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__36209\,
            I => \PWMInstance2.periodCounterZ0Z_10\
        );

    \I__8486\ : Odrv4
    port map (
            O => \N__36206\,
            I => \PWMInstance2.periodCounterZ0Z_10\
        );

    \I__8485\ : CascadeMux
    port map (
            O => \N__36201\,
            I => \N__36197\
        );

    \I__8484\ : CascadeMux
    port map (
            O => \N__36200\,
            I => \N__36193\
        );

    \I__8483\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36190\
        );

    \I__8482\ : InMux
    port map (
            O => \N__36196\,
            I => \N__36187\
        );

    \I__8481\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36184\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__36190\,
            I => \N__36181\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__36187\,
            I => \PWMInstance2.periodCounterZ0Z_11\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__36184\,
            I => \PWMInstance2.periodCounterZ0Z_11\
        );

    \I__8477\ : Odrv4
    port map (
            O => \N__36181\,
            I => \PWMInstance2.periodCounterZ0Z_11\
        );

    \I__8476\ : InMux
    port map (
            O => \N__36174\,
            I => \N__36171\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__36171\,
            I => \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_1\
        );

    \I__8474\ : InMux
    port map (
            O => \N__36168\,
            I => \N__36161\
        );

    \I__8473\ : InMux
    port map (
            O => \N__36167\,
            I => \N__36154\
        );

    \I__8472\ : InMux
    port map (
            O => \N__36166\,
            I => \N__36151\
        );

    \I__8471\ : InMux
    port map (
            O => \N__36165\,
            I => \N__36146\
        );

    \I__8470\ : CascadeMux
    port map (
            O => \N__36164\,
            I => \N__36143\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__36161\,
            I => \N__36139\
        );

    \I__8468\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36136\
        );

    \I__8467\ : InMux
    port map (
            O => \N__36159\,
            I => \N__36130\
        );

    \I__8466\ : InMux
    port map (
            O => \N__36158\,
            I => \N__36127\
        );

    \I__8465\ : InMux
    port map (
            O => \N__36157\,
            I => \N__36124\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__36154\,
            I => \N__36121\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__36151\,
            I => \N__36118\
        );

    \I__8462\ : InMux
    port map (
            O => \N__36150\,
            I => \N__36115\
        );

    \I__8461\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36112\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__36146\,
            I => \N__36109\
        );

    \I__8459\ : InMux
    port map (
            O => \N__36143\,
            I => \N__36106\
        );

    \I__8458\ : InMux
    port map (
            O => \N__36142\,
            I => \N__36103\
        );

    \I__8457\ : Span4Mux_v
    port map (
            O => \N__36139\,
            I => \N__36098\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__36136\,
            I => \N__36098\
        );

    \I__8455\ : InMux
    port map (
            O => \N__36135\,
            I => \N__36095\
        );

    \I__8454\ : InMux
    port map (
            O => \N__36134\,
            I => \N__36090\
        );

    \I__8453\ : InMux
    port map (
            O => \N__36133\,
            I => \N__36090\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__36130\,
            I => \N__36084\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__36127\,
            I => \N__36084\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__36124\,
            I => \N__36081\
        );

    \I__8449\ : Span4Mux_v
    port map (
            O => \N__36121\,
            I => \N__36076\
        );

    \I__8448\ : Span4Mux_v
    port map (
            O => \N__36118\,
            I => \N__36076\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36073\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__36112\,
            I => \N__36070\
        );

    \I__8445\ : Sp12to4
    port map (
            O => \N__36109\,
            I => \N__36065\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__36106\,
            I => \N__36065\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__36103\,
            I => \N__36062\
        );

    \I__8442\ : Span4Mux_h
    port map (
            O => \N__36098\,
            I => \N__36055\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__36095\,
            I => \N__36055\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__36090\,
            I => \N__36055\
        );

    \I__8439\ : InMux
    port map (
            O => \N__36089\,
            I => \N__36052\
        );

    \I__8438\ : Span4Mux_v
    port map (
            O => \N__36084\,
            I => \N__36049\
        );

    \I__8437\ : Span4Mux_h
    port map (
            O => \N__36081\,
            I => \N__36046\
        );

    \I__8436\ : Sp12to4
    port map (
            O => \N__36076\,
            I => \N__36037\
        );

    \I__8435\ : Span12Mux_s9_v
    port map (
            O => \N__36073\,
            I => \N__36037\
        );

    \I__8434\ : Span12Mux_s6_h
    port map (
            O => \N__36070\,
            I => \N__36037\
        );

    \I__8433\ : Span12Mux_s10_v
    port map (
            O => \N__36065\,
            I => \N__36037\
        );

    \I__8432\ : Span4Mux_h
    port map (
            O => \N__36062\,
            I => \N__36030\
        );

    \I__8431\ : Span4Mux_h
    port map (
            O => \N__36055\,
            I => \N__36030\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__36052\,
            I => \N__36030\
        );

    \I__8429\ : Odrv4
    port map (
            O => \N__36049\,
            I => \dataWriteZ0Z_10\
        );

    \I__8428\ : Odrv4
    port map (
            O => \N__36046\,
            I => \dataWriteZ0Z_10\
        );

    \I__8427\ : Odrv12
    port map (
            O => \N__36037\,
            I => \dataWriteZ0Z_10\
        );

    \I__8426\ : Odrv4
    port map (
            O => \N__36030\,
            I => \dataWriteZ0Z_10\
        );

    \I__8425\ : InMux
    port map (
            O => \N__36021\,
            I => \N__36018\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__36018\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_10\
        );

    \I__8423\ : CascadeMux
    port map (
            O => \N__36015\,
            I => \N__36007\
        );

    \I__8422\ : InMux
    port map (
            O => \N__36014\,
            I => \N__35999\
        );

    \I__8421\ : InMux
    port map (
            O => \N__36013\,
            I => \N__35995\
        );

    \I__8420\ : InMux
    port map (
            O => \N__36012\,
            I => \N__35990\
        );

    \I__8419\ : InMux
    port map (
            O => \N__36011\,
            I => \N__35987\
        );

    \I__8418\ : InMux
    port map (
            O => \N__36010\,
            I => \N__35978\
        );

    \I__8417\ : InMux
    port map (
            O => \N__36007\,
            I => \N__35978\
        );

    \I__8416\ : InMux
    port map (
            O => \N__36006\,
            I => \N__35978\
        );

    \I__8415\ : InMux
    port map (
            O => \N__36005\,
            I => \N__35978\
        );

    \I__8414\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35975\
        );

    \I__8413\ : InMux
    port map (
            O => \N__36003\,
            I => \N__35970\
        );

    \I__8412\ : InMux
    port map (
            O => \N__36002\,
            I => \N__35967\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__35999\,
            I => \N__35964\
        );

    \I__8410\ : InMux
    port map (
            O => \N__35998\,
            I => \N__35961\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__35995\,
            I => \N__35958\
        );

    \I__8408\ : InMux
    port map (
            O => \N__35994\,
            I => \N__35955\
        );

    \I__8407\ : InMux
    port map (
            O => \N__35993\,
            I => \N__35952\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__35990\,
            I => \N__35949\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__35987\,
            I => \N__35944\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__35978\,
            I => \N__35944\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__35975\,
            I => \N__35941\
        );

    \I__8402\ : InMux
    port map (
            O => \N__35974\,
            I => \N__35938\
        );

    \I__8401\ : CascadeMux
    port map (
            O => \N__35973\,
            I => \N__35935\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__35970\,
            I => \N__35930\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__35967\,
            I => \N__35930\
        );

    \I__8398\ : Span4Mux_v
    port map (
            O => \N__35964\,
            I => \N__35927\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__35961\,
            I => \N__35924\
        );

    \I__8396\ : Span4Mux_h
    port map (
            O => \N__35958\,
            I => \N__35919\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__35955\,
            I => \N__35919\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__35952\,
            I => \N__35916\
        );

    \I__8393\ : Span4Mux_v
    port map (
            O => \N__35949\,
            I => \N__35911\
        );

    \I__8392\ : Span4Mux_h
    port map (
            O => \N__35944\,
            I => \N__35911\
        );

    \I__8391\ : Span4Mux_h
    port map (
            O => \N__35941\,
            I => \N__35906\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__35938\,
            I => \N__35906\
        );

    \I__8389\ : InMux
    port map (
            O => \N__35935\,
            I => \N__35903\
        );

    \I__8388\ : Span12Mux_s10_v
    port map (
            O => \N__35930\,
            I => \N__35900\
        );

    \I__8387\ : Span4Mux_v
    port map (
            O => \N__35927\,
            I => \N__35897\
        );

    \I__8386\ : Span4Mux_h
    port map (
            O => \N__35924\,
            I => \N__35892\
        );

    \I__8385\ : Span4Mux_h
    port map (
            O => \N__35919\,
            I => \N__35892\
        );

    \I__8384\ : Span4Mux_v
    port map (
            O => \N__35916\,
            I => \N__35887\
        );

    \I__8383\ : Span4Mux_h
    port map (
            O => \N__35911\,
            I => \N__35887\
        );

    \I__8382\ : Span4Mux_h
    port map (
            O => \N__35906\,
            I => \N__35882\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__35903\,
            I => \N__35882\
        );

    \I__8380\ : Odrv12
    port map (
            O => \N__35900\,
            I => \dataWriteZ0Z_11\
        );

    \I__8379\ : Odrv4
    port map (
            O => \N__35897\,
            I => \dataWriteZ0Z_11\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__35892\,
            I => \dataWriteZ0Z_11\
        );

    \I__8377\ : Odrv4
    port map (
            O => \N__35887\,
            I => \dataWriteZ0Z_11\
        );

    \I__8376\ : Odrv4
    port map (
            O => \N__35882\,
            I => \dataWriteZ0Z_11\
        );

    \I__8375\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35868\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__35868\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_11\
        );

    \I__8373\ : CEMux
    port map (
            O => \N__35865\,
            I => \N__35862\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__35862\,
            I => \N__35858\
        );

    \I__8371\ : CEMux
    port map (
            O => \N__35861\,
            I => \N__35855\
        );

    \I__8370\ : Span4Mux_v
    port map (
            O => \N__35858\,
            I => \N__35848\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__35855\,
            I => \N__35848\
        );

    \I__8368\ : CEMux
    port map (
            O => \N__35854\,
            I => \N__35845\
        );

    \I__8367\ : CEMux
    port map (
            O => \N__35853\,
            I => \N__35842\
        );

    \I__8366\ : Span4Mux_h
    port map (
            O => \N__35848\,
            I => \N__35839\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__35845\,
            I => \PWMInstance2.pwmWrite_0_2\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__35842\,
            I => \PWMInstance2.pwmWrite_0_2\
        );

    \I__8363\ : Odrv4
    port map (
            O => \N__35839\,
            I => \PWMInstance2.pwmWrite_0_2\
        );

    \I__8362\ : InMux
    port map (
            O => \N__35832\,
            I => \N__35821\
        );

    \I__8361\ : InMux
    port map (
            O => \N__35831\,
            I => \N__35818\
        );

    \I__8360\ : InMux
    port map (
            O => \N__35830\,
            I => \N__35815\
        );

    \I__8359\ : InMux
    port map (
            O => \N__35829\,
            I => \N__35812\
        );

    \I__8358\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35809\
        );

    \I__8357\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35806\
        );

    \I__8356\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35803\
        );

    \I__8355\ : InMux
    port map (
            O => \N__35825\,
            I => \N__35800\
        );

    \I__8354\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35797\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__35821\,
            I => \N__35790\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__35818\,
            I => \N__35778\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__35815\,
            I => \N__35766\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__35812\,
            I => \N__35760\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__35809\,
            I => \N__35749\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__35806\,
            I => \N__35744\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__35803\,
            I => \N__35730\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__35800\,
            I => \N__35710\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__35797\,
            I => \N__35686\
        );

    \I__8344\ : SRMux
    port map (
            O => \N__35796\,
            I => \N__35469\
        );

    \I__8343\ : SRMux
    port map (
            O => \N__35795\,
            I => \N__35469\
        );

    \I__8342\ : SRMux
    port map (
            O => \N__35794\,
            I => \N__35469\
        );

    \I__8341\ : SRMux
    port map (
            O => \N__35793\,
            I => \N__35469\
        );

    \I__8340\ : Glb2LocalMux
    port map (
            O => \N__35790\,
            I => \N__35469\
        );

    \I__8339\ : SRMux
    port map (
            O => \N__35789\,
            I => \N__35469\
        );

    \I__8338\ : SRMux
    port map (
            O => \N__35788\,
            I => \N__35469\
        );

    \I__8337\ : SRMux
    port map (
            O => \N__35787\,
            I => \N__35469\
        );

    \I__8336\ : SRMux
    port map (
            O => \N__35786\,
            I => \N__35469\
        );

    \I__8335\ : SRMux
    port map (
            O => \N__35785\,
            I => \N__35469\
        );

    \I__8334\ : SRMux
    port map (
            O => \N__35784\,
            I => \N__35469\
        );

    \I__8333\ : SRMux
    port map (
            O => \N__35783\,
            I => \N__35469\
        );

    \I__8332\ : SRMux
    port map (
            O => \N__35782\,
            I => \N__35469\
        );

    \I__8331\ : SRMux
    port map (
            O => \N__35781\,
            I => \N__35469\
        );

    \I__8330\ : Glb2LocalMux
    port map (
            O => \N__35778\,
            I => \N__35469\
        );

    \I__8329\ : SRMux
    port map (
            O => \N__35777\,
            I => \N__35469\
        );

    \I__8328\ : SRMux
    port map (
            O => \N__35776\,
            I => \N__35469\
        );

    \I__8327\ : SRMux
    port map (
            O => \N__35775\,
            I => \N__35469\
        );

    \I__8326\ : SRMux
    port map (
            O => \N__35774\,
            I => \N__35469\
        );

    \I__8325\ : SRMux
    port map (
            O => \N__35773\,
            I => \N__35469\
        );

    \I__8324\ : SRMux
    port map (
            O => \N__35772\,
            I => \N__35469\
        );

    \I__8323\ : SRMux
    port map (
            O => \N__35771\,
            I => \N__35469\
        );

    \I__8322\ : SRMux
    port map (
            O => \N__35770\,
            I => \N__35469\
        );

    \I__8321\ : SRMux
    port map (
            O => \N__35769\,
            I => \N__35469\
        );

    \I__8320\ : Glb2LocalMux
    port map (
            O => \N__35766\,
            I => \N__35469\
        );

    \I__8319\ : SRMux
    port map (
            O => \N__35765\,
            I => \N__35469\
        );

    \I__8318\ : SRMux
    port map (
            O => \N__35764\,
            I => \N__35469\
        );

    \I__8317\ : SRMux
    port map (
            O => \N__35763\,
            I => \N__35469\
        );

    \I__8316\ : Glb2LocalMux
    port map (
            O => \N__35760\,
            I => \N__35469\
        );

    \I__8315\ : SRMux
    port map (
            O => \N__35759\,
            I => \N__35469\
        );

    \I__8314\ : SRMux
    port map (
            O => \N__35758\,
            I => \N__35469\
        );

    \I__8313\ : SRMux
    port map (
            O => \N__35757\,
            I => \N__35469\
        );

    \I__8312\ : SRMux
    port map (
            O => \N__35756\,
            I => \N__35469\
        );

    \I__8311\ : SRMux
    port map (
            O => \N__35755\,
            I => \N__35469\
        );

    \I__8310\ : SRMux
    port map (
            O => \N__35754\,
            I => \N__35469\
        );

    \I__8309\ : SRMux
    port map (
            O => \N__35753\,
            I => \N__35469\
        );

    \I__8308\ : SRMux
    port map (
            O => \N__35752\,
            I => \N__35469\
        );

    \I__8307\ : Glb2LocalMux
    port map (
            O => \N__35749\,
            I => \N__35469\
        );

    \I__8306\ : SRMux
    port map (
            O => \N__35748\,
            I => \N__35469\
        );

    \I__8305\ : SRMux
    port map (
            O => \N__35747\,
            I => \N__35469\
        );

    \I__8304\ : Glb2LocalMux
    port map (
            O => \N__35744\,
            I => \N__35469\
        );

    \I__8303\ : SRMux
    port map (
            O => \N__35743\,
            I => \N__35469\
        );

    \I__8302\ : SRMux
    port map (
            O => \N__35742\,
            I => \N__35469\
        );

    \I__8301\ : SRMux
    port map (
            O => \N__35741\,
            I => \N__35469\
        );

    \I__8300\ : SRMux
    port map (
            O => \N__35740\,
            I => \N__35469\
        );

    \I__8299\ : SRMux
    port map (
            O => \N__35739\,
            I => \N__35469\
        );

    \I__8298\ : SRMux
    port map (
            O => \N__35738\,
            I => \N__35469\
        );

    \I__8297\ : SRMux
    port map (
            O => \N__35737\,
            I => \N__35469\
        );

    \I__8296\ : SRMux
    port map (
            O => \N__35736\,
            I => \N__35469\
        );

    \I__8295\ : SRMux
    port map (
            O => \N__35735\,
            I => \N__35469\
        );

    \I__8294\ : SRMux
    port map (
            O => \N__35734\,
            I => \N__35469\
        );

    \I__8293\ : SRMux
    port map (
            O => \N__35733\,
            I => \N__35469\
        );

    \I__8292\ : Glb2LocalMux
    port map (
            O => \N__35730\,
            I => \N__35469\
        );

    \I__8291\ : SRMux
    port map (
            O => \N__35729\,
            I => \N__35469\
        );

    \I__8290\ : SRMux
    port map (
            O => \N__35728\,
            I => \N__35469\
        );

    \I__8289\ : SRMux
    port map (
            O => \N__35727\,
            I => \N__35469\
        );

    \I__8288\ : SRMux
    port map (
            O => \N__35726\,
            I => \N__35469\
        );

    \I__8287\ : SRMux
    port map (
            O => \N__35725\,
            I => \N__35469\
        );

    \I__8286\ : SRMux
    port map (
            O => \N__35724\,
            I => \N__35469\
        );

    \I__8285\ : SRMux
    port map (
            O => \N__35723\,
            I => \N__35469\
        );

    \I__8284\ : SRMux
    port map (
            O => \N__35722\,
            I => \N__35469\
        );

    \I__8283\ : SRMux
    port map (
            O => \N__35721\,
            I => \N__35469\
        );

    \I__8282\ : SRMux
    port map (
            O => \N__35720\,
            I => \N__35469\
        );

    \I__8281\ : SRMux
    port map (
            O => \N__35719\,
            I => \N__35469\
        );

    \I__8280\ : SRMux
    port map (
            O => \N__35718\,
            I => \N__35469\
        );

    \I__8279\ : SRMux
    port map (
            O => \N__35717\,
            I => \N__35469\
        );

    \I__8278\ : SRMux
    port map (
            O => \N__35716\,
            I => \N__35469\
        );

    \I__8277\ : SRMux
    port map (
            O => \N__35715\,
            I => \N__35469\
        );

    \I__8276\ : SRMux
    port map (
            O => \N__35714\,
            I => \N__35469\
        );

    \I__8275\ : SRMux
    port map (
            O => \N__35713\,
            I => \N__35469\
        );

    \I__8274\ : Glb2LocalMux
    port map (
            O => \N__35710\,
            I => \N__35469\
        );

    \I__8273\ : SRMux
    port map (
            O => \N__35709\,
            I => \N__35469\
        );

    \I__8272\ : SRMux
    port map (
            O => \N__35708\,
            I => \N__35469\
        );

    \I__8271\ : SRMux
    port map (
            O => \N__35707\,
            I => \N__35469\
        );

    \I__8270\ : SRMux
    port map (
            O => \N__35706\,
            I => \N__35469\
        );

    \I__8269\ : SRMux
    port map (
            O => \N__35705\,
            I => \N__35469\
        );

    \I__8268\ : SRMux
    port map (
            O => \N__35704\,
            I => \N__35469\
        );

    \I__8267\ : SRMux
    port map (
            O => \N__35703\,
            I => \N__35469\
        );

    \I__8266\ : SRMux
    port map (
            O => \N__35702\,
            I => \N__35469\
        );

    \I__8265\ : SRMux
    port map (
            O => \N__35701\,
            I => \N__35469\
        );

    \I__8264\ : SRMux
    port map (
            O => \N__35700\,
            I => \N__35469\
        );

    \I__8263\ : SRMux
    port map (
            O => \N__35699\,
            I => \N__35469\
        );

    \I__8262\ : SRMux
    port map (
            O => \N__35698\,
            I => \N__35469\
        );

    \I__8261\ : SRMux
    port map (
            O => \N__35697\,
            I => \N__35469\
        );

    \I__8260\ : SRMux
    port map (
            O => \N__35696\,
            I => \N__35469\
        );

    \I__8259\ : SRMux
    port map (
            O => \N__35695\,
            I => \N__35469\
        );

    \I__8258\ : SRMux
    port map (
            O => \N__35694\,
            I => \N__35469\
        );

    \I__8257\ : SRMux
    port map (
            O => \N__35693\,
            I => \N__35469\
        );

    \I__8256\ : SRMux
    port map (
            O => \N__35692\,
            I => \N__35469\
        );

    \I__8255\ : SRMux
    port map (
            O => \N__35691\,
            I => \N__35469\
        );

    \I__8254\ : SRMux
    port map (
            O => \N__35690\,
            I => \N__35469\
        );

    \I__8253\ : SRMux
    port map (
            O => \N__35689\,
            I => \N__35469\
        );

    \I__8252\ : Glb2LocalMux
    port map (
            O => \N__35686\,
            I => \N__35469\
        );

    \I__8251\ : SRMux
    port map (
            O => \N__35685\,
            I => \N__35469\
        );

    \I__8250\ : SRMux
    port map (
            O => \N__35684\,
            I => \N__35469\
        );

    \I__8249\ : SRMux
    port map (
            O => \N__35683\,
            I => \N__35469\
        );

    \I__8248\ : SRMux
    port map (
            O => \N__35682\,
            I => \N__35469\
        );

    \I__8247\ : SRMux
    port map (
            O => \N__35681\,
            I => \N__35469\
        );

    \I__8246\ : SRMux
    port map (
            O => \N__35680\,
            I => \N__35469\
        );

    \I__8245\ : SRMux
    port map (
            O => \N__35679\,
            I => \N__35469\
        );

    \I__8244\ : SRMux
    port map (
            O => \N__35678\,
            I => \N__35469\
        );

    \I__8243\ : SRMux
    port map (
            O => \N__35677\,
            I => \N__35469\
        );

    \I__8242\ : SRMux
    port map (
            O => \N__35676\,
            I => \N__35469\
        );

    \I__8241\ : GlobalMux
    port map (
            O => \N__35469\,
            I => \N__35466\
        );

    \I__8240\ : gio2CtrlBuf
    port map (
            O => \N__35466\,
            I => \RST_c_i_g\
        );

    \I__8239\ : IoInMux
    port map (
            O => \N__35463\,
            I => \N__35460\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__35460\,
            I => \PWM2_obufLegalizeSB_DFFNet\
        );

    \I__8237\ : InMux
    port map (
            O => \N__35457\,
            I => \N__35452\
        );

    \I__8236\ : InMux
    port map (
            O => \N__35456\,
            I => \N__35449\
        );

    \I__8235\ : InMux
    port map (
            O => \N__35455\,
            I => \N__35446\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__35452\,
            I => \PWMInstance2.periodCounterZ0Z_9\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__35449\,
            I => \PWMInstance2.periodCounterZ0Z_9\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__35446\,
            I => \PWMInstance2.periodCounterZ0Z_9\
        );

    \I__8231\ : InMux
    port map (
            O => \N__35439\,
            I => \PWMInstance2.un1_periodCounter_2_cry_8\
        );

    \I__8230\ : InMux
    port map (
            O => \N__35436\,
            I => \PWMInstance2.un1_periodCounter_2_cry_9\
        );

    \I__8229\ : InMux
    port map (
            O => \N__35433\,
            I => \PWMInstance2.un1_periodCounter_2_cry_10\
        );

    \I__8228\ : InMux
    port map (
            O => \N__35430\,
            I => \PWMInstance2.un1_periodCounter_2_cry_11\
        );

    \I__8227\ : CascadeMux
    port map (
            O => \N__35427\,
            I => \N__35423\
        );

    \I__8226\ : InMux
    port map (
            O => \N__35426\,
            I => \N__35419\
        );

    \I__8225\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35416\
        );

    \I__8224\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35413\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__35419\,
            I => \PWMInstance2.periodCounterZ0Z_13\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__35416\,
            I => \PWMInstance2.periodCounterZ0Z_13\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__35413\,
            I => \PWMInstance2.periodCounterZ0Z_13\
        );

    \I__8220\ : InMux
    port map (
            O => \N__35406\,
            I => \PWMInstance2.un1_periodCounter_2_cry_12\
        );

    \I__8219\ : InMux
    port map (
            O => \N__35403\,
            I => \PWMInstance2.un1_periodCounter_2_cry_13\
        );

    \I__8218\ : CascadeMux
    port map (
            O => \N__35400\,
            I => \N__35396\
        );

    \I__8217\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35392\
        );

    \I__8216\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35389\
        );

    \I__8215\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35386\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__35392\,
            I => \PWMInstance2.periodCounterZ0Z_15\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__35389\,
            I => \PWMInstance2.periodCounterZ0Z_15\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__35386\,
            I => \PWMInstance2.periodCounterZ0Z_15\
        );

    \I__8211\ : InMux
    port map (
            O => \N__35379\,
            I => \PWMInstance2.un1_periodCounter_2_cry_14\
        );

    \I__8210\ : CascadeMux
    port map (
            O => \N__35376\,
            I => \N__35373\
        );

    \I__8209\ : InMux
    port map (
            O => \N__35373\,
            I => \N__35365\
        );

    \I__8208\ : InMux
    port map (
            O => \N__35372\,
            I => \N__35362\
        );

    \I__8207\ : InMux
    port map (
            O => \N__35371\,
            I => \N__35359\
        );

    \I__8206\ : InMux
    port map (
            O => \N__35370\,
            I => \N__35354\
        );

    \I__8205\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35354\
        );

    \I__8204\ : InMux
    port map (
            O => \N__35368\,
            I => \N__35351\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__35365\,
            I => \N__35348\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__35362\,
            I => \PWMInstance2.out_0_sqmuxa\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__35359\,
            I => \PWMInstance2.out_0_sqmuxa\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__35354\,
            I => \PWMInstance2.out_0_sqmuxa\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__35351\,
            I => \PWMInstance2.out_0_sqmuxa\
        );

    \I__8198\ : Odrv4
    port map (
            O => \N__35348\,
            I => \PWMInstance2.out_0_sqmuxa\
        );

    \I__8197\ : InMux
    port map (
            O => \N__35337\,
            I => \bfn_18_13_0_\
        );

    \I__8196\ : CascadeMux
    port map (
            O => \N__35334\,
            I => \N__35330\
        );

    \I__8195\ : InMux
    port map (
            O => \N__35333\,
            I => \N__35326\
        );

    \I__8194\ : InMux
    port map (
            O => \N__35330\,
            I => \N__35321\
        );

    \I__8193\ : InMux
    port map (
            O => \N__35329\,
            I => \N__35321\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__35326\,
            I => \PWMInstance2.periodCounterZ0Z_16\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__35321\,
            I => \PWMInstance2.periodCounterZ0Z_16\
        );

    \I__8190\ : SRMux
    port map (
            O => \N__35316\,
            I => \N__35244\
        );

    \I__8189\ : SRMux
    port map (
            O => \N__35315\,
            I => \N__35244\
        );

    \I__8188\ : SRMux
    port map (
            O => \N__35314\,
            I => \N__35244\
        );

    \I__8187\ : SRMux
    port map (
            O => \N__35313\,
            I => \N__35244\
        );

    \I__8186\ : SRMux
    port map (
            O => \N__35312\,
            I => \N__35244\
        );

    \I__8185\ : SRMux
    port map (
            O => \N__35311\,
            I => \N__35244\
        );

    \I__8184\ : SRMux
    port map (
            O => \N__35310\,
            I => \N__35244\
        );

    \I__8183\ : SRMux
    port map (
            O => \N__35309\,
            I => \N__35244\
        );

    \I__8182\ : SRMux
    port map (
            O => \N__35308\,
            I => \N__35244\
        );

    \I__8181\ : SRMux
    port map (
            O => \N__35307\,
            I => \N__35244\
        );

    \I__8180\ : SRMux
    port map (
            O => \N__35306\,
            I => \N__35244\
        );

    \I__8179\ : SRMux
    port map (
            O => \N__35305\,
            I => \N__35244\
        );

    \I__8178\ : SRMux
    port map (
            O => \N__35304\,
            I => \N__35244\
        );

    \I__8177\ : SRMux
    port map (
            O => \N__35303\,
            I => \N__35244\
        );

    \I__8176\ : SRMux
    port map (
            O => \N__35302\,
            I => \N__35244\
        );

    \I__8175\ : SRMux
    port map (
            O => \N__35301\,
            I => \N__35244\
        );

    \I__8174\ : SRMux
    port map (
            O => \N__35300\,
            I => \N__35244\
        );

    \I__8173\ : SRMux
    port map (
            O => \N__35299\,
            I => \N__35244\
        );

    \I__8172\ : SRMux
    port map (
            O => \N__35298\,
            I => \N__35244\
        );

    \I__8171\ : SRMux
    port map (
            O => \N__35297\,
            I => \N__35244\
        );

    \I__8170\ : SRMux
    port map (
            O => \N__35296\,
            I => \N__35244\
        );

    \I__8169\ : SRMux
    port map (
            O => \N__35295\,
            I => \N__35244\
        );

    \I__8168\ : SRMux
    port map (
            O => \N__35294\,
            I => \N__35244\
        );

    \I__8167\ : SRMux
    port map (
            O => \N__35293\,
            I => \N__35244\
        );

    \I__8166\ : GlobalMux
    port map (
            O => \N__35244\,
            I => \N__35241\
        );

    \I__8165\ : gio2CtrlBuf
    port map (
            O => \N__35241\,
            I => \PWMInstance0_N_42_g\
        );

    \I__8164\ : CascadeMux
    port map (
            O => \N__35238\,
            I => \N__35234\
        );

    \I__8163\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35230\
        );

    \I__8162\ : InMux
    port map (
            O => \N__35234\,
            I => \N__35227\
        );

    \I__8161\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35224\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__35230\,
            I => \N__35219\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__35227\,
            I => \N__35219\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__35224\,
            I => \PWMInstance2.periodCounterZ0Z_5\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__35219\,
            I => \PWMInstance2.periodCounterZ0Z_5\
        );

    \I__8156\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__35211\,
            I => \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_1\
        );

    \I__8154\ : CascadeMux
    port map (
            O => \N__35208\,
            I => \N__35203\
        );

    \I__8153\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35200\
        );

    \I__8152\ : InMux
    port map (
            O => \N__35206\,
            I => \N__35197\
        );

    \I__8151\ : InMux
    port map (
            O => \N__35203\,
            I => \N__35194\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__35200\,
            I => \PWMInstance2.periodCounterZ0Z_1\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__35197\,
            I => \PWMInstance2.periodCounterZ0Z_1\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__35194\,
            I => \PWMInstance2.periodCounterZ0Z_1\
        );

    \I__8147\ : InMux
    port map (
            O => \N__35187\,
            I => \PWMInstance2.un1_periodCounter_2_cry_0\
        );

    \I__8146\ : InMux
    port map (
            O => \N__35184\,
            I => \PWMInstance2.un1_periodCounter_2_cry_1\
        );

    \I__8145\ : InMux
    port map (
            O => \N__35181\,
            I => \N__35174\
        );

    \I__8144\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35174\
        );

    \I__8143\ : InMux
    port map (
            O => \N__35179\,
            I => \N__35171\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__35174\,
            I => \N__35168\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__35171\,
            I => \PWMInstance2.periodCounterZ0Z_3\
        );

    \I__8140\ : Odrv4
    port map (
            O => \N__35168\,
            I => \PWMInstance2.periodCounterZ0Z_3\
        );

    \I__8139\ : InMux
    port map (
            O => \N__35163\,
            I => \PWMInstance2.un1_periodCounter_2_cry_2\
        );

    \I__8138\ : InMux
    port map (
            O => \N__35160\,
            I => \PWMInstance2.un1_periodCounter_2_cry_3\
        );

    \I__8137\ : InMux
    port map (
            O => \N__35157\,
            I => \PWMInstance2.un1_periodCounter_2_cry_4\
        );

    \I__8136\ : CascadeMux
    port map (
            O => \N__35154\,
            I => \N__35149\
        );

    \I__8135\ : CascadeMux
    port map (
            O => \N__35153\,
            I => \N__35146\
        );

    \I__8134\ : InMux
    port map (
            O => \N__35152\,
            I => \N__35143\
        );

    \I__8133\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35138\
        );

    \I__8132\ : InMux
    port map (
            O => \N__35146\,
            I => \N__35138\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__35143\,
            I => \PWMInstance2.periodCounterZ0Z_6\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__35138\,
            I => \PWMInstance2.periodCounterZ0Z_6\
        );

    \I__8129\ : InMux
    port map (
            O => \N__35133\,
            I => \PWMInstance2.un1_periodCounter_2_cry_5\
        );

    \I__8128\ : InMux
    port map (
            O => \N__35130\,
            I => \N__35125\
        );

    \I__8127\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35122\
        );

    \I__8126\ : InMux
    port map (
            O => \N__35128\,
            I => \N__35119\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__35125\,
            I => \PWMInstance2.periodCounterZ0Z_7\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__35122\,
            I => \PWMInstance2.periodCounterZ0Z_7\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__35119\,
            I => \PWMInstance2.periodCounterZ0Z_7\
        );

    \I__8122\ : InMux
    port map (
            O => \N__35112\,
            I => \PWMInstance2.un1_periodCounter_2_cry_6\
        );

    \I__8121\ : CascadeMux
    port map (
            O => \N__35109\,
            I => \N__35104\
        );

    \I__8120\ : InMux
    port map (
            O => \N__35108\,
            I => \N__35101\
        );

    \I__8119\ : InMux
    port map (
            O => \N__35107\,
            I => \N__35096\
        );

    \I__8118\ : InMux
    port map (
            O => \N__35104\,
            I => \N__35096\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__35101\,
            I => \PWMInstance2.periodCounterZ0Z_8\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__35096\,
            I => \PWMInstance2.periodCounterZ0Z_8\
        );

    \I__8115\ : InMux
    port map (
            O => \N__35091\,
            I => \bfn_18_12_0_\
        );

    \I__8114\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35076\
        );

    \I__8113\ : InMux
    port map (
            O => \N__35087\,
            I => \N__35076\
        );

    \I__8112\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35076\
        );

    \I__8111\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35076\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__35076\,
            I => \N__35073\
        );

    \I__8109\ : Span4Mux_v
    port map (
            O => \N__35073\,
            I => \N__35070\
        );

    \I__8108\ : Span4Mux_h
    port map (
            O => \N__35070\,
            I => \N__35067\
        );

    \I__8107\ : Span4Mux_h
    port map (
            O => \N__35067\,
            I => \N__35064\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__35064\,
            I => \MOSIrZ0Z_1\
        );

    \I__8105\ : InMux
    port map (
            O => \N__35061\,
            I => \N__35057\
        );

    \I__8104\ : InMux
    port map (
            O => \N__35060\,
            I => \N__35054\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__35057\,
            I => \N__35051\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__35054\,
            I => \N__35047\
        );

    \I__8101\ : Span4Mux_v
    port map (
            O => \N__35051\,
            I => \N__35044\
        );

    \I__8100\ : InMux
    port map (
            O => \N__35050\,
            I => \N__35041\
        );

    \I__8099\ : Span4Mux_h
    port map (
            O => \N__35047\,
            I => \N__35038\
        );

    \I__8098\ : Span4Mux_v
    port map (
            O => \N__35044\,
            I => \N__35033\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__35041\,
            I => \N__35033\
        );

    \I__8096\ : Span4Mux_h
    port map (
            O => \N__35038\,
            I => \N__35030\
        );

    \I__8095\ : Odrv4
    port map (
            O => \N__35033\,
            I => \dataRead1_10\
        );

    \I__8094\ : Odrv4
    port map (
            O => \N__35030\,
            I => \dataRead1_10\
        );

    \I__8093\ : CascadeMux
    port map (
            O => \N__35025\,
            I => \N__35021\
        );

    \I__8092\ : CascadeMux
    port map (
            O => \N__35024\,
            I => \N__35018\
        );

    \I__8091\ : InMux
    port map (
            O => \N__35021\,
            I => \N__35015\
        );

    \I__8090\ : InMux
    port map (
            O => \N__35018\,
            I => \N__35012\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__35015\,
            I => \N__35009\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__35012\,
            I => \N__35005\
        );

    \I__8087\ : Span4Mux_v
    port map (
            O => \N__35009\,
            I => \N__35002\
        );

    \I__8086\ : InMux
    port map (
            O => \N__35008\,
            I => \N__34999\
        );

    \I__8085\ : Span4Mux_v
    port map (
            O => \N__35005\,
            I => \N__34994\
        );

    \I__8084\ : Span4Mux_h
    port map (
            O => \N__35002\,
            I => \N__34994\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__34999\,
            I => \dataRead5_10\
        );

    \I__8082\ : Odrv4
    port map (
            O => \N__34994\,
            I => \dataRead5_10\
        );

    \I__8081\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34986\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__34986\,
            I => \N__34983\
        );

    \I__8079\ : Odrv4
    port map (
            O => \N__34983\,
            I => \OutReg_0_5_i_m3_ns_1_10\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__34980\,
            I => \N__34975\
        );

    \I__8077\ : InMux
    port map (
            O => \N__34979\,
            I => \N__34972\
        );

    \I__8076\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34969\
        );

    \I__8075\ : InMux
    port map (
            O => \N__34975\,
            I => \N__34966\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__34972\,
            I => \N__34961\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34961\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__34966\,
            I => \N__34958\
        );

    \I__8071\ : Span4Mux_v
    port map (
            O => \N__34961\,
            I => \N__34953\
        );

    \I__8070\ : Span4Mux_h
    port map (
            O => \N__34958\,
            I => \N__34953\
        );

    \I__8069\ : Span4Mux_h
    port map (
            O => \N__34953\,
            I => \N__34950\
        );

    \I__8068\ : Odrv4
    port map (
            O => \N__34950\,
            I => \data_receivedZ0Z_4\
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__34947\,
            I => \un1_OutReg51_4_0_i_o3_2_cascade_\
        );

    \I__8066\ : InMux
    port map (
            O => \N__34944\,
            I => \N__34941\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__34941\,
            I => \OutReg_21_m_0_a2_1_0\
        );

    \I__8064\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34935\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__34935\,
            I => \OutReg_esr_RNO_2Z0Z_10\
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__34932\,
            I => \N__34929\
        );

    \I__8061\ : InMux
    port map (
            O => \N__34929\,
            I => \N__34926\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__34926\,
            I => \N__34923\
        );

    \I__8059\ : Span4Mux_h
    port map (
            O => \N__34923\,
            I => \N__34920\
        );

    \I__8058\ : Odrv4
    port map (
            O => \N__34920\,
            I => \OutRegZ0Z_9\
        );

    \I__8057\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34914\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__34914\,
            I => \OutReg_esr_RNO_0Z0Z_10\
        );

    \I__8055\ : InMux
    port map (
            O => \N__34911\,
            I => \N__34908\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__34908\,
            I => \N__34905\
        );

    \I__8053\ : Span4Mux_h
    port map (
            O => \N__34905\,
            I => \N__34902\
        );

    \I__8052\ : Span4Mux_h
    port map (
            O => \N__34902\,
            I => \N__34899\
        );

    \I__8051\ : Odrv4
    port map (
            O => \N__34899\,
            I => \OutRegZ0Z_10\
        );

    \I__8050\ : CascadeMux
    port map (
            O => \N__34896\,
            I => \N__34890\
        );

    \I__8049\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34886\
        );

    \I__8048\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34880\
        );

    \I__8047\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34877\
        );

    \I__8046\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34874\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__34889\,
            I => \N__34871\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__34886\,
            I => \N__34867\
        );

    \I__8043\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34864\
        );

    \I__8042\ : CascadeMux
    port map (
            O => \N__34884\,
            I => \N__34859\
        );

    \I__8041\ : InMux
    port map (
            O => \N__34883\,
            I => \N__34856\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__34880\,
            I => \N__34851\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__34877\,
            I => \N__34851\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__34874\,
            I => \N__34848\
        );

    \I__8037\ : InMux
    port map (
            O => \N__34871\,
            I => \N__34845\
        );

    \I__8036\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34842\
        );

    \I__8035\ : Span4Mux_v
    port map (
            O => \N__34867\,
            I => \N__34839\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__34864\,
            I => \N__34836\
        );

    \I__8033\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34833\
        );

    \I__8032\ : InMux
    port map (
            O => \N__34862\,
            I => \N__34828\
        );

    \I__8031\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34828\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__34856\,
            I => \N__34823\
        );

    \I__8029\ : Span4Mux_h
    port map (
            O => \N__34851\,
            I => \N__34823\
        );

    \I__8028\ : Span4Mux_h
    port map (
            O => \N__34848\,
            I => \N__34818\
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__34845\,
            I => \N__34818\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__34842\,
            I => \data_received_fastZ0Z_2\
        );

    \I__8025\ : Odrv4
    port map (
            O => \N__34839\,
            I => \data_received_fastZ0Z_2\
        );

    \I__8024\ : Odrv12
    port map (
            O => \N__34836\,
            I => \data_received_fastZ0Z_2\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__34833\,
            I => \data_received_fastZ0Z_2\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__34828\,
            I => \data_received_fastZ0Z_2\
        );

    \I__8021\ : Odrv4
    port map (
            O => \N__34823\,
            I => \data_received_fastZ0Z_2\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__34818\,
            I => \data_received_fastZ0Z_2\
        );

    \I__8019\ : InMux
    port map (
            O => \N__34803\,
            I => \N__34799\
        );

    \I__8018\ : InMux
    port map (
            O => \N__34802\,
            I => \N__34796\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__34799\,
            I => \N__34793\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__34796\,
            I => \N__34790\
        );

    \I__8015\ : Span4Mux_h
    port map (
            O => \N__34793\,
            I => \N__34784\
        );

    \I__8014\ : Span4Mux_h
    port map (
            O => \N__34790\,
            I => \N__34784\
        );

    \I__8013\ : InMux
    port map (
            O => \N__34789\,
            I => \N__34781\
        );

    \I__8012\ : Span4Mux_h
    port map (
            O => \N__34784\,
            I => \N__34778\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__34781\,
            I => \dataRead3_10\
        );

    \I__8010\ : Odrv4
    port map (
            O => \N__34778\,
            I => \dataRead3_10\
        );

    \I__8009\ : CascadeMux
    port map (
            O => \N__34773\,
            I => \N__34768\
        );

    \I__8008\ : CascadeMux
    port map (
            O => \N__34772\,
            I => \N__34765\
        );

    \I__8007\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34758\
        );

    \I__8006\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34755\
        );

    \I__8005\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34752\
        );

    \I__8004\ : InMux
    port map (
            O => \N__34764\,
            I => \N__34749\
        );

    \I__8003\ : InMux
    port map (
            O => \N__34763\,
            I => \N__34746\
        );

    \I__8002\ : InMux
    port map (
            O => \N__34762\,
            I => \N__34743\
        );

    \I__8001\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34739\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__34758\,
            I => \N__34734\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__34755\,
            I => \N__34734\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__34752\,
            I => \N__34728\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__34749\,
            I => \N__34725\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__34746\,
            I => \N__34722\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__34743\,
            I => \N__34719\
        );

    \I__7994\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34716\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__34739\,
            I => \N__34711\
        );

    \I__7992\ : Span4Mux_h
    port map (
            O => \N__34734\,
            I => \N__34711\
        );

    \I__7991\ : InMux
    port map (
            O => \N__34733\,
            I => \N__34706\
        );

    \I__7990\ : InMux
    port map (
            O => \N__34732\,
            I => \N__34706\
        );

    \I__7989\ : InMux
    port map (
            O => \N__34731\,
            I => \N__34703\
        );

    \I__7988\ : Span4Mux_v
    port map (
            O => \N__34728\,
            I => \N__34696\
        );

    \I__7987\ : Span4Mux_v
    port map (
            O => \N__34725\,
            I => \N__34696\
        );

    \I__7986\ : Span4Mux_v
    port map (
            O => \N__34722\,
            I => \N__34696\
        );

    \I__7985\ : Odrv4
    port map (
            O => \N__34719\,
            I => \data_received_fastZ0Z_0\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__34716\,
            I => \data_received_fastZ0Z_0\
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__34711\,
            I => \data_received_fastZ0Z_0\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__34706\,
            I => \data_received_fastZ0Z_0\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__34703\,
            I => \data_received_fastZ0Z_0\
        );

    \I__7980\ : Odrv4
    port map (
            O => \N__34696\,
            I => \data_received_fastZ0Z_0\
        );

    \I__7979\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34680\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__34680\,
            I => \N__34677\
        );

    \I__7977\ : Span4Mux_v
    port map (
            O => \N__34677\,
            I => \N__34672\
        );

    \I__7976\ : InMux
    port map (
            O => \N__34676\,
            I => \N__34669\
        );

    \I__7975\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34666\
        );

    \I__7974\ : Span4Mux_h
    port map (
            O => \N__34672\,
            I => \N__34663\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__34669\,
            I => \N__34660\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__34666\,
            I => \N__34655\
        );

    \I__7971\ : Span4Mux_h
    port map (
            O => \N__34663\,
            I => \N__34655\
        );

    \I__7970\ : Odrv4
    port map (
            O => \N__34660\,
            I => \dataRead2_10\
        );

    \I__7969\ : Odrv4
    port map (
            O => \N__34655\,
            I => \dataRead2_10\
        );

    \I__7968\ : InMux
    port map (
            O => \N__34650\,
            I => \N__34646\
        );

    \I__7967\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34642\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__34646\,
            I => \N__34639\
        );

    \I__7965\ : InMux
    port map (
            O => \N__34645\,
            I => \N__34636\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__34642\,
            I => \N__34633\
        );

    \I__7963\ : Span4Mux_v
    port map (
            O => \N__34639\,
            I => \N__34628\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__34636\,
            I => \N__34628\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__34633\,
            I => \N__34625\
        );

    \I__7960\ : Span4Mux_h
    port map (
            O => \N__34628\,
            I => \N__34622\
        );

    \I__7959\ : Span4Mux_h
    port map (
            O => \N__34625\,
            I => \N__34619\
        );

    \I__7958\ : Odrv4
    port map (
            O => \N__34622\,
            I => \dataRead7_10\
        );

    \I__7957\ : Odrv4
    port map (
            O => \N__34619\,
            I => \dataRead7_10\
        );

    \I__7956\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34611\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__34611\,
            I => \N__34606\
        );

    \I__7954\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34603\
        );

    \I__7953\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34600\
        );

    \I__7952\ : Span4Mux_h
    port map (
            O => \N__34606\,
            I => \N__34597\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__34603\,
            I => \N__34594\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__34600\,
            I => \N__34591\
        );

    \I__7949\ : Span4Mux_h
    port map (
            O => \N__34597\,
            I => \N__34588\
        );

    \I__7948\ : Odrv4
    port map (
            O => \N__34594\,
            I => \dataRead6_10\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__34591\,
            I => \dataRead6_10\
        );

    \I__7946\ : Odrv4
    port map (
            O => \N__34588\,
            I => \dataRead6_10\
        );

    \I__7945\ : CascadeMux
    port map (
            O => \N__34581\,
            I => \OutReg_0_4_i_m3_ns_1_10_cascade_\
        );

    \I__7944\ : InMux
    port map (
            O => \N__34578\,
            I => \N__34575\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__34575\,
            I => \OutReg_esr_RNO_1Z0Z_10\
        );

    \I__7942\ : CascadeMux
    port map (
            O => \N__34572\,
            I => \N__34568\
        );

    \I__7941\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34564\
        );

    \I__7940\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34561\
        );

    \I__7939\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34558\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__34564\,
            I => \PWMInstance2.periodCounter12\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__34561\,
            I => \PWMInstance2.periodCounter12\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__34558\,
            I => \PWMInstance2.periodCounter12\
        );

    \I__7935\ : InMux
    port map (
            O => \N__34551\,
            I => \N__34546\
        );

    \I__7934\ : InMux
    port map (
            O => \N__34550\,
            I => \N__34541\
        );

    \I__7933\ : InMux
    port map (
            O => \N__34549\,
            I => \N__34541\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__34546\,
            I => \PWMInstance2.periodCounterZ0Z_0\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__34541\,
            I => \PWMInstance2.periodCounterZ0Z_0\
        );

    \I__7930\ : CascadeMux
    port map (
            O => \N__34536\,
            I => \N__34531\
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__34535\,
            I => \N__34528\
        );

    \I__7928\ : InMux
    port map (
            O => \N__34534\,
            I => \N__34525\
        );

    \I__7927\ : InMux
    port map (
            O => \N__34531\,
            I => \N__34520\
        );

    \I__7926\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34520\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__34525\,
            I => \QuadInstance0.delayedCh_AZ0Z_1\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__34520\,
            I => \QuadInstance0.delayedCh_AZ0Z_1\
        );

    \I__7923\ : InMux
    port map (
            O => \N__34515\,
            I => \N__34512\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__34512\,
            I => \N__34508\
        );

    \I__7921\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34505\
        );

    \I__7920\ : Span4Mux_h
    port map (
            O => \N__34508\,
            I => \N__34502\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34497\
        );

    \I__7918\ : Span4Mux_v
    port map (
            O => \N__34502\,
            I => \N__34492\
        );

    \I__7917\ : InMux
    port map (
            O => \N__34501\,
            I => \N__34489\
        );

    \I__7916\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34486\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__34497\,
            I => \N__34483\
        );

    \I__7914\ : InMux
    port map (
            O => \N__34496\,
            I => \N__34480\
        );

    \I__7913\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34477\
        );

    \I__7912\ : Span4Mux_v
    port map (
            O => \N__34492\,
            I => \N__34472\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__34489\,
            I => \N__34472\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__34486\,
            I => \N__34466\
        );

    \I__7909\ : Sp12to4
    port map (
            O => \N__34483\,
            I => \N__34459\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__34480\,
            I => \N__34459\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__34477\,
            I => \N__34459\
        );

    \I__7906\ : Span4Mux_v
    port map (
            O => \N__34472\,
            I => \N__34456\
        );

    \I__7905\ : InMux
    port map (
            O => \N__34471\,
            I => \N__34453\
        );

    \I__7904\ : InMux
    port map (
            O => \N__34470\,
            I => \N__34450\
        );

    \I__7903\ : InMux
    port map (
            O => \N__34469\,
            I => \N__34447\
        );

    \I__7902\ : Span12Mux_h
    port map (
            O => \N__34466\,
            I => \N__34442\
        );

    \I__7901\ : Span12Mux_h
    port map (
            O => \N__34459\,
            I => \N__34442\
        );

    \I__7900\ : Span4Mux_v
    port map (
            O => \N__34456\,
            I => \N__34439\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__34453\,
            I => \N__34432\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__34450\,
            I => \N__34432\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__34447\,
            I => \N__34432\
        );

    \I__7896\ : Span12Mux_v
    port map (
            O => \N__34442\,
            I => \N__34429\
        );

    \I__7895\ : IoSpan4Mux
    port map (
            O => \N__34439\,
            I => \N__34426\
        );

    \I__7894\ : Span12Mux_h
    port map (
            O => \N__34432\,
            I => \N__34423\
        );

    \I__7893\ : Odrv12
    port map (
            O => \N__34429\,
            I => \RST_c\
        );

    \I__7892\ : Odrv4
    port map (
            O => \N__34426\,
            I => \RST_c\
        );

    \I__7891\ : Odrv12
    port map (
            O => \N__34423\,
            I => \RST_c\
        );

    \I__7890\ : InMux
    port map (
            O => \N__34416\,
            I => \N__34410\
        );

    \I__7889\ : InMux
    port map (
            O => \N__34415\,
            I => \N__34407\
        );

    \I__7888\ : InMux
    port map (
            O => \N__34414\,
            I => \N__34404\
        );

    \I__7887\ : InMux
    port map (
            O => \N__34413\,
            I => \N__34396\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__34410\,
            I => \N__34391\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__34407\,
            I => \N__34388\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__34404\,
            I => \N__34385\
        );

    \I__7883\ : InMux
    port map (
            O => \N__34403\,
            I => \N__34382\
        );

    \I__7882\ : InMux
    port map (
            O => \N__34402\,
            I => \N__34379\
        );

    \I__7881\ : InMux
    port map (
            O => \N__34401\,
            I => \N__34375\
        );

    \I__7880\ : InMux
    port map (
            O => \N__34400\,
            I => \N__34370\
        );

    \I__7879\ : InMux
    port map (
            O => \N__34399\,
            I => \N__34367\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__34396\,
            I => \N__34362\
        );

    \I__7877\ : InMux
    port map (
            O => \N__34395\,
            I => \N__34359\
        );

    \I__7876\ : InMux
    port map (
            O => \N__34394\,
            I => \N__34356\
        );

    \I__7875\ : Span4Mux_v
    port map (
            O => \N__34391\,
            I => \N__34351\
        );

    \I__7874\ : Span4Mux_h
    port map (
            O => \N__34388\,
            I => \N__34351\
        );

    \I__7873\ : Span4Mux_h
    port map (
            O => \N__34385\,
            I => \N__34346\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__34382\,
            I => \N__34346\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__34379\,
            I => \N__34343\
        );

    \I__7870\ : InMux
    port map (
            O => \N__34378\,
            I => \N__34340\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__34375\,
            I => \N__34337\
        );

    \I__7868\ : InMux
    port map (
            O => \N__34374\,
            I => \N__34332\
        );

    \I__7867\ : InMux
    port map (
            O => \N__34373\,
            I => \N__34332\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__34370\,
            I => \N__34329\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__34367\,
            I => \N__34326\
        );

    \I__7864\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34323\
        );

    \I__7863\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34320\
        );

    \I__7862\ : Span4Mux_v
    port map (
            O => \N__34362\,
            I => \N__34317\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__34359\,
            I => \N__34312\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__34356\,
            I => \N__34312\
        );

    \I__7859\ : Span4Mux_v
    port map (
            O => \N__34351\,
            I => \N__34309\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__34346\,
            I => \N__34304\
        );

    \I__7857\ : Span4Mux_h
    port map (
            O => \N__34343\,
            I => \N__34304\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__34340\,
            I => \N__34301\
        );

    \I__7855\ : Span4Mux_v
    port map (
            O => \N__34337\,
            I => \N__34298\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__34332\,
            I => \N__34295\
        );

    \I__7853\ : Span4Mux_h
    port map (
            O => \N__34329\,
            I => \N__34292\
        );

    \I__7852\ : Span4Mux_h
    port map (
            O => \N__34326\,
            I => \N__34285\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__34323\,
            I => \N__34285\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__34320\,
            I => \N__34285\
        );

    \I__7849\ : Span4Mux_h
    port map (
            O => \N__34317\,
            I => \N__34276\
        );

    \I__7848\ : Span4Mux_v
    port map (
            O => \N__34312\,
            I => \N__34276\
        );

    \I__7847\ : Span4Mux_h
    port map (
            O => \N__34309\,
            I => \N__34276\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__34304\,
            I => \N__34276\
        );

    \I__7845\ : Span4Mux_h
    port map (
            O => \N__34301\,
            I => \N__34269\
        );

    \I__7844\ : Span4Mux_h
    port map (
            O => \N__34298\,
            I => \N__34269\
        );

    \I__7843\ : Span4Mux_v
    port map (
            O => \N__34295\,
            I => \N__34269\
        );

    \I__7842\ : Span4Mux_h
    port map (
            O => \N__34292\,
            I => \N__34264\
        );

    \I__7841\ : Span4Mux_h
    port map (
            O => \N__34285\,
            I => \N__34264\
        );

    \I__7840\ : Odrv4
    port map (
            O => \N__34276\,
            I => \dataWriteZ0Z_14\
        );

    \I__7839\ : Odrv4
    port map (
            O => \N__34269\,
            I => \dataWriteZ0Z_14\
        );

    \I__7838\ : Odrv4
    port map (
            O => \N__34264\,
            I => \dataWriteZ0Z_14\
        );

    \I__7837\ : InMux
    port map (
            O => \N__34257\,
            I => \N__34254\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__34254\,
            I => \QuadInstance0.Quad_RNO_0_0_14\
        );

    \I__7835\ : InMux
    port map (
            O => \N__34251\,
            I => \N__34246\
        );

    \I__7834\ : CascadeMux
    port map (
            O => \N__34250\,
            I => \N__34243\
        );

    \I__7833\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34240\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__34246\,
            I => \N__34237\
        );

    \I__7831\ : InMux
    port map (
            O => \N__34243\,
            I => \N__34234\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__34240\,
            I => \N__34229\
        );

    \I__7829\ : Span4Mux_v
    port map (
            O => \N__34237\,
            I => \N__34229\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__34234\,
            I => \dataRead0_14\
        );

    \I__7827\ : Odrv4
    port map (
            O => \N__34229\,
            I => \dataRead0_14\
        );

    \I__7826\ : InMux
    port map (
            O => \N__34224\,
            I => \N__34221\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__34221\,
            I => \QuadInstance0.Quad_RNI4P8Q1Z0Z_14\
        );

    \I__7824\ : CascadeMux
    port map (
            O => \N__34218\,
            I => \N__34214\
        );

    \I__7823\ : InMux
    port map (
            O => \N__34217\,
            I => \N__34211\
        );

    \I__7822\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34208\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__34211\,
            I => \N__34204\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__34208\,
            I => \N__34201\
        );

    \I__7819\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34198\
        );

    \I__7818\ : Span4Mux_h
    port map (
            O => \N__34204\,
            I => \N__34195\
        );

    \I__7817\ : Span4Mux_h
    port map (
            O => \N__34201\,
            I => \N__34192\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__34198\,
            I => \N__34189\
        );

    \I__7815\ : Span4Mux_h
    port map (
            O => \N__34195\,
            I => \N__34186\
        );

    \I__7814\ : Span4Mux_h
    port map (
            O => \N__34192\,
            I => \N__34183\
        );

    \I__7813\ : Odrv12
    port map (
            O => \N__34189\,
            I => \dataRead0_3\
        );

    \I__7812\ : Odrv4
    port map (
            O => \N__34186\,
            I => \dataRead0_3\
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__34183\,
            I => \dataRead0_3\
        );

    \I__7810\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34173\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__34173\,
            I => \QuadInstance0.Quad_RNIIGBH1Z0Z_3\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__34170\,
            I => \N__34167\
        );

    \I__7807\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34164\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__34164\,
            I => \N__34160\
        );

    \I__7805\ : InMux
    port map (
            O => \N__34163\,
            I => \N__34157\
        );

    \I__7804\ : Span4Mux_v
    port map (
            O => \N__34160\,
            I => \N__34154\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__34157\,
            I => \N__34150\
        );

    \I__7802\ : Sp12to4
    port map (
            O => \N__34154\,
            I => \N__34147\
        );

    \I__7801\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34144\
        );

    \I__7800\ : Span4Mux_v
    port map (
            O => \N__34150\,
            I => \N__34141\
        );

    \I__7799\ : Odrv12
    port map (
            O => \N__34147\,
            I => \dataRead0_4\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__34144\,
            I => \dataRead0_4\
        );

    \I__7797\ : Odrv4
    port map (
            O => \N__34141\,
            I => \dataRead0_4\
        );

    \I__7796\ : CascadeMux
    port map (
            O => \N__34134\,
            I => \N__34131\
        );

    \I__7795\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34128\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__34128\,
            I => \QuadInstance0.Quad_RNIJHBH1Z0Z_4\
        );

    \I__7793\ : InMux
    port map (
            O => \N__34125\,
            I => \N__34122\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__34122\,
            I => \N__34118\
        );

    \I__7791\ : InMux
    port map (
            O => \N__34121\,
            I => \N__34115\
        );

    \I__7790\ : Span4Mux_v
    port map (
            O => \N__34118\,
            I => \N__34111\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__34115\,
            I => \N__34108\
        );

    \I__7788\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34105\
        );

    \I__7787\ : Odrv4
    port map (
            O => \N__34111\,
            I => \dataRead0_5\
        );

    \I__7786\ : Odrv4
    port map (
            O => \N__34108\,
            I => \dataRead0_5\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__34105\,
            I => \dataRead0_5\
        );

    \I__7784\ : CascadeMux
    port map (
            O => \N__34098\,
            I => \N__34095\
        );

    \I__7783\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34092\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__34092\,
            I => \QuadInstance0.Quad_RNIKIBH1Z0Z_5\
        );

    \I__7781\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34082\
        );

    \I__7780\ : CascadeMux
    port map (
            O => \N__34088\,
            I => \N__34078\
        );

    \I__7779\ : CascadeMux
    port map (
            O => \N__34087\,
            I => \N__34074\
        );

    \I__7778\ : CascadeMux
    port map (
            O => \N__34086\,
            I => \N__34071\
        );

    \I__7777\ : CascadeMux
    port map (
            O => \N__34085\,
            I => \N__34068\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__34082\,
            I => \N__34065\
        );

    \I__7775\ : CascadeMux
    port map (
            O => \N__34081\,
            I => \N__34062\
        );

    \I__7774\ : InMux
    port map (
            O => \N__34078\,
            I => \N__34054\
        );

    \I__7773\ : InMux
    port map (
            O => \N__34077\,
            I => \N__34054\
        );

    \I__7772\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34054\
        );

    \I__7771\ : InMux
    port map (
            O => \N__34071\,
            I => \N__34049\
        );

    \I__7770\ : InMux
    port map (
            O => \N__34068\,
            I => \N__34049\
        );

    \I__7769\ : Span4Mux_v
    port map (
            O => \N__34065\,
            I => \N__34043\
        );

    \I__7768\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34038\
        );

    \I__7767\ : InMux
    port map (
            O => \N__34061\,
            I => \N__34038\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__34054\,
            I => \N__34033\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__34049\,
            I => \N__34033\
        );

    \I__7764\ : CascadeMux
    port map (
            O => \N__34048\,
            I => \N__34025\
        );

    \I__7763\ : InMux
    port map (
            O => \N__34047\,
            I => \N__34022\
        );

    \I__7762\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34019\
        );

    \I__7761\ : Span4Mux_h
    port map (
            O => \N__34043\,
            I => \N__34014\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__34038\,
            I => \N__34014\
        );

    \I__7759\ : Span4Mux_h
    port map (
            O => \N__34033\,
            I => \N__34011\
        );

    \I__7758\ : InMux
    port map (
            O => \N__34032\,
            I => \N__34002\
        );

    \I__7757\ : InMux
    port map (
            O => \N__34031\,
            I => \N__34002\
        );

    \I__7756\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34002\
        );

    \I__7755\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34002\
        );

    \I__7754\ : InMux
    port map (
            O => \N__34028\,
            I => \N__33997\
        );

    \I__7753\ : InMux
    port map (
            O => \N__34025\,
            I => \N__33997\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__34022\,
            I => \QuadInstance0.count_enable\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__34019\,
            I => \QuadInstance0.count_enable\
        );

    \I__7750\ : Odrv4
    port map (
            O => \N__34014\,
            I => \QuadInstance0.count_enable\
        );

    \I__7749\ : Odrv4
    port map (
            O => \N__34011\,
            I => \QuadInstance0.count_enable\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__34002\,
            I => \QuadInstance0.count_enable\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__33997\,
            I => \QuadInstance0.count_enable\
        );

    \I__7746\ : CascadeMux
    port map (
            O => \N__33984\,
            I => \N__33981\
        );

    \I__7745\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33977\
        );

    \I__7744\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33974\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__33977\,
            I => \N__33971\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__33974\,
            I => \N__33967\
        );

    \I__7741\ : Span4Mux_v
    port map (
            O => \N__33971\,
            I => \N__33964\
        );

    \I__7740\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33961\
        );

    \I__7739\ : Span4Mux_h
    port map (
            O => \N__33967\,
            I => \N__33958\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__33964\,
            I => \dataRead0_6\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__33961\,
            I => \dataRead0_6\
        );

    \I__7736\ : Odrv4
    port map (
            O => \N__33958\,
            I => \dataRead0_6\
        );

    \I__7735\ : CascadeMux
    port map (
            O => \N__33951\,
            I => \N__33946\
        );

    \I__7734\ : CascadeMux
    port map (
            O => \N__33950\,
            I => \N__33939\
        );

    \I__7733\ : InMux
    port map (
            O => \N__33949\,
            I => \N__33932\
        );

    \I__7732\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33932\
        );

    \I__7731\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33932\
        );

    \I__7730\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33927\
        );

    \I__7729\ : InMux
    port map (
            O => \N__33943\,
            I => \N__33927\
        );

    \I__7728\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33919\
        );

    \I__7727\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33919\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__33932\,
            I => \N__33914\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__33927\,
            I => \N__33914\
        );

    \I__7724\ : CascadeMux
    port map (
            O => \N__33926\,
            I => \N__33910\
        );

    \I__7723\ : CascadeMux
    port map (
            O => \N__33925\,
            I => \N__33906\
        );

    \I__7722\ : InMux
    port map (
            O => \N__33924\,
            I => \N__33900\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__33919\,
            I => \N__33897\
        );

    \I__7720\ : Span4Mux_h
    port map (
            O => \N__33914\,
            I => \N__33894\
        );

    \I__7719\ : InMux
    port map (
            O => \N__33913\,
            I => \N__33883\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33910\,
            I => \N__33883\
        );

    \I__7717\ : InMux
    port map (
            O => \N__33909\,
            I => \N__33883\
        );

    \I__7716\ : InMux
    port map (
            O => \N__33906\,
            I => \N__33883\
        );

    \I__7715\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33883\
        );

    \I__7714\ : InMux
    port map (
            O => \N__33904\,
            I => \N__33878\
        );

    \I__7713\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33878\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__33900\,
            I => \QuadInstance0.un1_count_enable_i_a2_0_1\
        );

    \I__7711\ : Odrv4
    port map (
            O => \N__33897\,
            I => \QuadInstance0.un1_count_enable_i_a2_0_1\
        );

    \I__7710\ : Odrv4
    port map (
            O => \N__33894\,
            I => \QuadInstance0.un1_count_enable_i_a2_0_1\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__33883\,
            I => \QuadInstance0.un1_count_enable_i_a2_0_1\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__33878\,
            I => \QuadInstance0.un1_count_enable_i_a2_0_1\
        );

    \I__7707\ : CascadeMux
    port map (
            O => \N__33867\,
            I => \N__33864\
        );

    \I__7706\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33861\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__33861\,
            I => \QuadInstance0.Quad_RNILJBH1Z0Z_6\
        );

    \I__7704\ : InMux
    port map (
            O => \N__33858\,
            I => \N__33852\
        );

    \I__7703\ : InMux
    port map (
            O => \N__33857\,
            I => \N__33843\
        );

    \I__7702\ : InMux
    port map (
            O => \N__33856\,
            I => \N__33837\
        );

    \I__7701\ : InMux
    port map (
            O => \N__33855\,
            I => \N__33837\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__33852\,
            I => \N__33834\
        );

    \I__7699\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33831\
        );

    \I__7698\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33823\
        );

    \I__7697\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33819\
        );

    \I__7696\ : InMux
    port map (
            O => \N__33848\,
            I => \N__33816\
        );

    \I__7695\ : InMux
    port map (
            O => \N__33847\,
            I => \N__33813\
        );

    \I__7694\ : InMux
    port map (
            O => \N__33846\,
            I => \N__33810\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__33843\,
            I => \N__33807\
        );

    \I__7692\ : InMux
    port map (
            O => \N__33842\,
            I => \N__33804\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__33837\,
            I => \N__33801\
        );

    \I__7690\ : Span4Mux_v
    port map (
            O => \N__33834\,
            I => \N__33796\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__33831\,
            I => \N__33796\
        );

    \I__7688\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33793\
        );

    \I__7687\ : InMux
    port map (
            O => \N__33829\,
            I => \N__33788\
        );

    \I__7686\ : InMux
    port map (
            O => \N__33828\,
            I => \N__33788\
        );

    \I__7685\ : InMux
    port map (
            O => \N__33827\,
            I => \N__33785\
        );

    \I__7684\ : InMux
    port map (
            O => \N__33826\,
            I => \N__33780\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__33823\,
            I => \N__33777\
        );

    \I__7682\ : InMux
    port map (
            O => \N__33822\,
            I => \N__33774\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__33819\,
            I => \N__33771\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__33816\,
            I => \N__33762\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__33813\,
            I => \N__33762\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__33810\,
            I => \N__33762\
        );

    \I__7677\ : Span4Mux_h
    port map (
            O => \N__33807\,
            I => \N__33762\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__33804\,
            I => \N__33752\
        );

    \I__7675\ : Span4Mux_v
    port map (
            O => \N__33801\,
            I => \N__33752\
        );

    \I__7674\ : Span4Mux_h
    port map (
            O => \N__33796\,
            I => \N__33752\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__33793\,
            I => \N__33744\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__33788\,
            I => \N__33744\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__33785\,
            I => \N__33741\
        );

    \I__7670\ : InMux
    port map (
            O => \N__33784\,
            I => \N__33736\
        );

    \I__7669\ : InMux
    port map (
            O => \N__33783\,
            I => \N__33736\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__33780\,
            I => \N__33733\
        );

    \I__7667\ : Span4Mux_v
    port map (
            O => \N__33777\,
            I => \N__33730\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__33774\,
            I => \N__33723\
        );

    \I__7665\ : Span4Mux_v
    port map (
            O => \N__33771\,
            I => \N__33723\
        );

    \I__7664\ : Span4Mux_v
    port map (
            O => \N__33762\,
            I => \N__33723\
        );

    \I__7663\ : InMux
    port map (
            O => \N__33761\,
            I => \N__33716\
        );

    \I__7662\ : InMux
    port map (
            O => \N__33760\,
            I => \N__33716\
        );

    \I__7661\ : InMux
    port map (
            O => \N__33759\,
            I => \N__33716\
        );

    \I__7660\ : Span4Mux_v
    port map (
            O => \N__33752\,
            I => \N__33713\
        );

    \I__7659\ : InMux
    port map (
            O => \N__33751\,
            I => \N__33708\
        );

    \I__7658\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33708\
        );

    \I__7657\ : InMux
    port map (
            O => \N__33749\,
            I => \N__33705\
        );

    \I__7656\ : Span4Mux_h
    port map (
            O => \N__33744\,
            I => \N__33702\
        );

    \I__7655\ : Span12Mux_s11_v
    port map (
            O => \N__33741\,
            I => \N__33699\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__33736\,
            I => \N__33690\
        );

    \I__7653\ : Span4Mux_v
    port map (
            O => \N__33733\,
            I => \N__33690\
        );

    \I__7652\ : Span4Mux_h
    port map (
            O => \N__33730\,
            I => \N__33690\
        );

    \I__7651\ : Span4Mux_h
    port map (
            O => \N__33723\,
            I => \N__33690\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__33716\,
            I => \N__33685\
        );

    \I__7649\ : Span4Mux_h
    port map (
            O => \N__33713\,
            I => \N__33685\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__33708\,
            I => \data_receivedZ0Z_21\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__33705\,
            I => \data_receivedZ0Z_21\
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__33702\,
            I => \data_receivedZ0Z_21\
        );

    \I__7645\ : Odrv12
    port map (
            O => \N__33699\,
            I => \data_receivedZ0Z_21\
        );

    \I__7644\ : Odrv4
    port map (
            O => \N__33690\,
            I => \data_receivedZ0Z_21\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__33685\,
            I => \data_receivedZ0Z_21\
        );

    \I__7642\ : InMux
    port map (
            O => \N__33672\,
            I => \N__33667\
        );

    \I__7641\ : CascadeMux
    port map (
            O => \N__33671\,
            I => \N__33663\
        );

    \I__7640\ : InMux
    port map (
            O => \N__33670\,
            I => \N__33653\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__33667\,
            I => \N__33648\
        );

    \I__7638\ : InMux
    port map (
            O => \N__33666\,
            I => \N__33645\
        );

    \I__7637\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33640\
        );

    \I__7636\ : InMux
    port map (
            O => \N__33662\,
            I => \N__33640\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__33661\,
            I => \N__33634\
        );

    \I__7634\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33631\
        );

    \I__7633\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33628\
        );

    \I__7632\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33623\
        );

    \I__7631\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33623\
        );

    \I__7630\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33620\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__33653\,
            I => \N__33616\
        );

    \I__7628\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33611\
        );

    \I__7627\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33611\
        );

    \I__7626\ : Span4Mux_v
    port map (
            O => \N__33648\,
            I => \N__33604\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__33645\,
            I => \N__33604\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__33640\,
            I => \N__33604\
        );

    \I__7623\ : InMux
    port map (
            O => \N__33639\,
            I => \N__33601\
        );

    \I__7622\ : CascadeMux
    port map (
            O => \N__33638\,
            I => \N__33596\
        );

    \I__7621\ : CascadeMux
    port map (
            O => \N__33637\,
            I => \N__33593\
        );

    \I__7620\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33590\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__33631\,
            I => \N__33587\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__33628\,
            I => \N__33583\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__33623\,
            I => \N__33578\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__33620\,
            I => \N__33578\
        );

    \I__7615\ : InMux
    port map (
            O => \N__33619\,
            I => \N__33575\
        );

    \I__7614\ : Span4Mux_v
    port map (
            O => \N__33616\,
            I => \N__33572\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__33611\,
            I => \N__33565\
        );

    \I__7612\ : Span4Mux_v
    port map (
            O => \N__33604\,
            I => \N__33565\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__33601\,
            I => \N__33565\
        );

    \I__7610\ : CascadeMux
    port map (
            O => \N__33600\,
            I => \N__33562\
        );

    \I__7609\ : InMux
    port map (
            O => \N__33599\,
            I => \N__33554\
        );

    \I__7608\ : InMux
    port map (
            O => \N__33596\,
            I => \N__33549\
        );

    \I__7607\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33549\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__33590\,
            I => \N__33546\
        );

    \I__7605\ : Span4Mux_v
    port map (
            O => \N__33587\,
            I => \N__33543\
        );

    \I__7604\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33540\
        );

    \I__7603\ : Span4Mux_v
    port map (
            O => \N__33583\,
            I => \N__33537\
        );

    \I__7602\ : Span4Mux_v
    port map (
            O => \N__33578\,
            I => \N__33534\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__33575\,
            I => \N__33531\
        );

    \I__7600\ : Span4Mux_h
    port map (
            O => \N__33572\,
            I => \N__33526\
        );

    \I__7599\ : Span4Mux_v
    port map (
            O => \N__33565\,
            I => \N__33526\
        );

    \I__7598\ : InMux
    port map (
            O => \N__33562\,
            I => \N__33521\
        );

    \I__7597\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33521\
        );

    \I__7596\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33518\
        );

    \I__7595\ : InMux
    port map (
            O => \N__33559\,
            I => \N__33511\
        );

    \I__7594\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33511\
        );

    \I__7593\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33511\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__33554\,
            I => \N__33508\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__33549\,
            I => \N__33503\
        );

    \I__7590\ : Span4Mux_h
    port map (
            O => \N__33546\,
            I => \N__33503\
        );

    \I__7589\ : Span4Mux_h
    port map (
            O => \N__33543\,
            I => \N__33500\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__33540\,
            I => \N__33493\
        );

    \I__7587\ : Span4Mux_h
    port map (
            O => \N__33537\,
            I => \N__33493\
        );

    \I__7586\ : Span4Mux_v
    port map (
            O => \N__33534\,
            I => \N__33493\
        );

    \I__7585\ : Span12Mux_s11_v
    port map (
            O => \N__33531\,
            I => \N__33490\
        );

    \I__7584\ : Span4Mux_h
    port map (
            O => \N__33526\,
            I => \N__33487\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__33521\,
            I => \data_receivedZ0Z_20\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__33518\,
            I => \data_receivedZ0Z_20\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__33511\,
            I => \data_receivedZ0Z_20\
        );

    \I__7580\ : Odrv4
    port map (
            O => \N__33508\,
            I => \data_receivedZ0Z_20\
        );

    \I__7579\ : Odrv4
    port map (
            O => \N__33503\,
            I => \data_receivedZ0Z_20\
        );

    \I__7578\ : Odrv4
    port map (
            O => \N__33500\,
            I => \data_receivedZ0Z_20\
        );

    \I__7577\ : Odrv4
    port map (
            O => \N__33493\,
            I => \data_receivedZ0Z_20\
        );

    \I__7576\ : Odrv12
    port map (
            O => \N__33490\,
            I => \data_receivedZ0Z_20\
        );

    \I__7575\ : Odrv4
    port map (
            O => \N__33487\,
            I => \data_receivedZ0Z_20\
        );

    \I__7574\ : CascadeMux
    port map (
            O => \N__33468\,
            I => \N__33460\
        );

    \I__7573\ : CascadeMux
    port map (
            O => \N__33467\,
            I => \N__33453\
        );

    \I__7572\ : CascadeMux
    port map (
            O => \N__33466\,
            I => \N__33443\
        );

    \I__7571\ : CascadeMux
    port map (
            O => \N__33465\,
            I => \N__33437\
        );

    \I__7570\ : CascadeMux
    port map (
            O => \N__33464\,
            I => \N__33433\
        );

    \I__7569\ : CascadeMux
    port map (
            O => \N__33463\,
            I => \N__33429\
        );

    \I__7568\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33426\
        );

    \I__7567\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33421\
        );

    \I__7566\ : InMux
    port map (
            O => \N__33458\,
            I => \N__33421\
        );

    \I__7565\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33416\
        );

    \I__7564\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33416\
        );

    \I__7563\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33413\
        );

    \I__7562\ : CascadeMux
    port map (
            O => \N__33452\,
            I => \N__33410\
        );

    \I__7561\ : CascadeMux
    port map (
            O => \N__33451\,
            I => \N__33407\
        );

    \I__7560\ : CascadeMux
    port map (
            O => \N__33450\,
            I => \N__33404\
        );

    \I__7559\ : CascadeMux
    port map (
            O => \N__33449\,
            I => \N__33401\
        );

    \I__7558\ : CascadeMux
    port map (
            O => \N__33448\,
            I => \N__33397\
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__33447\,
            I => \N__33394\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__33446\,
            I => \N__33391\
        );

    \I__7555\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33388\
        );

    \I__7554\ : CascadeMux
    port map (
            O => \N__33442\,
            I => \N__33385\
        );

    \I__7553\ : CascadeMux
    port map (
            O => \N__33441\,
            I => \N__33382\
        );

    \I__7552\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33377\
        );

    \I__7551\ : InMux
    port map (
            O => \N__33437\,
            I => \N__33377\
        );

    \I__7550\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33374\
        );

    \I__7549\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33371\
        );

    \I__7548\ : CascadeMux
    port map (
            O => \N__33432\,
            I => \N__33368\
        );

    \I__7547\ : InMux
    port map (
            O => \N__33429\,
            I => \N__33364\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__33426\,
            I => \N__33357\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__33421\,
            I => \N__33357\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__33416\,
            I => \N__33357\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__33413\,
            I => \N__33354\
        );

    \I__7542\ : InMux
    port map (
            O => \N__33410\,
            I => \N__33351\
        );

    \I__7541\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33346\
        );

    \I__7540\ : InMux
    port map (
            O => \N__33404\,
            I => \N__33346\
        );

    \I__7539\ : InMux
    port map (
            O => \N__33401\,
            I => \N__33343\
        );

    \I__7538\ : CascadeMux
    port map (
            O => \N__33400\,
            I => \N__33340\
        );

    \I__7537\ : InMux
    port map (
            O => \N__33397\,
            I => \N__33337\
        );

    \I__7536\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33332\
        );

    \I__7535\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33332\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__33388\,
            I => \N__33329\
        );

    \I__7533\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33326\
        );

    \I__7532\ : InMux
    port map (
            O => \N__33382\,
            I => \N__33323\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__33377\,
            I => \N__33316\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__33374\,
            I => \N__33316\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__33371\,
            I => \N__33316\
        );

    \I__7528\ : InMux
    port map (
            O => \N__33368\,
            I => \N__33311\
        );

    \I__7527\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33311\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__33364\,
            I => \N__33304\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__33357\,
            I => \N__33304\
        );

    \I__7524\ : Span4Mux_v
    port map (
            O => \N__33354\,
            I => \N__33304\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__33351\,
            I => \N__33301\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__33346\,
            I => \N__33298\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__33343\,
            I => \N__33295\
        );

    \I__7520\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33292\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__33337\,
            I => \N__33287\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__33332\,
            I => \N__33287\
        );

    \I__7517\ : Span4Mux_h
    port map (
            O => \N__33329\,
            I => \N__33284\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__33326\,
            I => \N__33276\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__33323\,
            I => \N__33276\
        );

    \I__7514\ : Span4Mux_v
    port map (
            O => \N__33316\,
            I => \N__33276\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__33311\,
            I => \N__33267\
        );

    \I__7512\ : Span4Mux_h
    port map (
            O => \N__33304\,
            I => \N__33267\
        );

    \I__7511\ : Span4Mux_v
    port map (
            O => \N__33301\,
            I => \N__33267\
        );

    \I__7510\ : Span4Mux_v
    port map (
            O => \N__33298\,
            I => \N__33267\
        );

    \I__7509\ : Sp12to4
    port map (
            O => \N__33295\,
            I => \N__33264\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__33292\,
            I => \N__33259\
        );

    \I__7507\ : Span4Mux_h
    port map (
            O => \N__33287\,
            I => \N__33259\
        );

    \I__7506\ : Span4Mux_v
    port map (
            O => \N__33284\,
            I => \N__33256\
        );

    \I__7505\ : InMux
    port map (
            O => \N__33283\,
            I => \N__33253\
        );

    \I__7504\ : Sp12to4
    port map (
            O => \N__33276\,
            I => \N__33246\
        );

    \I__7503\ : Sp12to4
    port map (
            O => \N__33267\,
            I => \N__33246\
        );

    \I__7502\ : Span12Mux_s9_v
    port map (
            O => \N__33264\,
            I => \N__33246\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__33259\,
            I => \N__33241\
        );

    \I__7500\ : Span4Mux_h
    port map (
            O => \N__33256\,
            I => \N__33241\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__33253\,
            I => \data_receivedZ0Z_22\
        );

    \I__7498\ : Odrv12
    port map (
            O => \N__33246\,
            I => \data_receivedZ0Z_22\
        );

    \I__7497\ : Odrv4
    port map (
            O => \N__33241\,
            I => \data_receivedZ0Z_22\
        );

    \I__7496\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33226\
        );

    \I__7495\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33226\
        );

    \I__7494\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33221\
        );

    \I__7493\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33218\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__33226\,
            I => \N__33215\
        );

    \I__7491\ : InMux
    port map (
            O => \N__33225\,
            I => \N__33211\
        );

    \I__7490\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33208\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__33221\,
            I => \N__33204\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__33218\,
            I => \N__33200\
        );

    \I__7487\ : Span4Mux_h
    port map (
            O => \N__33215\,
            I => \N__33197\
        );

    \I__7486\ : InMux
    port map (
            O => \N__33214\,
            I => \N__33194\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__33211\,
            I => \N__33189\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__33208\,
            I => \N__33186\
        );

    \I__7483\ : InMux
    port map (
            O => \N__33207\,
            I => \N__33183\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__33204\,
            I => \N__33180\
        );

    \I__7481\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33177\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__33200\,
            I => \N__33174\
        );

    \I__7479\ : Span4Mux_v
    port map (
            O => \N__33197\,
            I => \N__33169\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33169\
        );

    \I__7477\ : InMux
    port map (
            O => \N__33193\,
            I => \N__33164\
        );

    \I__7476\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33164\
        );

    \I__7475\ : Span4Mux_v
    port map (
            O => \N__33189\,
            I => \N__33157\
        );

    \I__7474\ : Span4Mux_v
    port map (
            O => \N__33186\,
            I => \N__33157\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__33183\,
            I => \N__33157\
        );

    \I__7472\ : Span4Mux_h
    port map (
            O => \N__33180\,
            I => \N__33154\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__33177\,
            I => \N__33151\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__33174\,
            I => \N__33144\
        );

    \I__7469\ : Span4Mux_h
    port map (
            O => \N__33169\,
            I => \N__33144\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__33164\,
            I => \N__33144\
        );

    \I__7467\ : Span4Mux_h
    port map (
            O => \N__33157\,
            I => \N__33141\
        );

    \I__7466\ : Odrv4
    port map (
            O => \N__33154\,
            I => \data_received_esr_RNIMIH31_0Z0Z_19\
        );

    \I__7465\ : Odrv4
    port map (
            O => \N__33151\,
            I => \data_received_esr_RNIMIH31_0Z0Z_19\
        );

    \I__7464\ : Odrv4
    port map (
            O => \N__33144\,
            I => \data_received_esr_RNIMIH31_0Z0Z_19\
        );

    \I__7463\ : Odrv4
    port map (
            O => \N__33141\,
            I => \data_received_esr_RNIMIH31_0Z0Z_19\
        );

    \I__7462\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33121\
        );

    \I__7461\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33121\
        );

    \I__7460\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33117\
        );

    \I__7459\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33104\
        );

    \I__7458\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33104\
        );

    \I__7457\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33097\
        );

    \I__7456\ : InMux
    port map (
            O => \N__33126\,
            I => \N__33094\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__33121\,
            I => \N__33091\
        );

    \I__7454\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33088\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33085\
        );

    \I__7452\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33074\
        );

    \I__7451\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33074\
        );

    \I__7450\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33074\
        );

    \I__7449\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33074\
        );

    \I__7448\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33074\
        );

    \I__7447\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33069\
        );

    \I__7446\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33069\
        );

    \I__7445\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33066\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__33104\,
            I => \N__33063\
        );

    \I__7443\ : InMux
    port map (
            O => \N__33103\,
            I => \N__33054\
        );

    \I__7442\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33054\
        );

    \I__7441\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33054\
        );

    \I__7440\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33054\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__33097\,
            I => \N__33049\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__33094\,
            I => \N__33039\
        );

    \I__7437\ : Span4Mux_v
    port map (
            O => \N__33091\,
            I => \N__33039\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__33088\,
            I => \N__33030\
        );

    \I__7435\ : Span4Mux_h
    port map (
            O => \N__33085\,
            I => \N__33030\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__33074\,
            I => \N__33030\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__33069\,
            I => \N__33030\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__33066\,
            I => \N__33027\
        );

    \I__7431\ : Span4Mux_v
    port map (
            O => \N__33063\,
            I => \N__33022\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__33054\,
            I => \N__33022\
        );

    \I__7429\ : CascadeMux
    port map (
            O => \N__33053\,
            I => \N__33019\
        );

    \I__7428\ : CascadeMux
    port map (
            O => \N__33052\,
            I => \N__33016\
        );

    \I__7427\ : Span4Mux_h
    port map (
            O => \N__33049\,
            I => \N__33009\
        );

    \I__7426\ : InMux
    port map (
            O => \N__33048\,
            I => \N__33000\
        );

    \I__7425\ : InMux
    port map (
            O => \N__33047\,
            I => \N__33000\
        );

    \I__7424\ : InMux
    port map (
            O => \N__33046\,
            I => \N__33000\
        );

    \I__7423\ : InMux
    port map (
            O => \N__33045\,
            I => \N__33000\
        );

    \I__7422\ : InMux
    port map (
            O => \N__33044\,
            I => \N__32997\
        );

    \I__7421\ : Span4Mux_h
    port map (
            O => \N__33039\,
            I => \N__32992\
        );

    \I__7420\ : Span4Mux_v
    port map (
            O => \N__33030\,
            I => \N__32992\
        );

    \I__7419\ : Span4Mux_v
    port map (
            O => \N__33027\,
            I => \N__32987\
        );

    \I__7418\ : Span4Mux_h
    port map (
            O => \N__33022\,
            I => \N__32987\
        );

    \I__7417\ : InMux
    port map (
            O => \N__33019\,
            I => \N__32974\
        );

    \I__7416\ : InMux
    port map (
            O => \N__33016\,
            I => \N__32974\
        );

    \I__7415\ : InMux
    port map (
            O => \N__33015\,
            I => \N__32974\
        );

    \I__7414\ : InMux
    port map (
            O => \N__33014\,
            I => \N__32974\
        );

    \I__7413\ : InMux
    port map (
            O => \N__33013\,
            I => \N__32974\
        );

    \I__7412\ : InMux
    port map (
            O => \N__33012\,
            I => \N__32974\
        );

    \I__7411\ : Span4Mux_h
    port map (
            O => \N__33009\,
            I => \N__32969\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__33000\,
            I => \N__32969\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__32997\,
            I => \quadWriteZ0Z_0\
        );

    \I__7408\ : Odrv4
    port map (
            O => \N__32992\,
            I => \quadWriteZ0Z_0\
        );

    \I__7407\ : Odrv4
    port map (
            O => \N__32987\,
            I => \quadWriteZ0Z_0\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__32974\,
            I => \quadWriteZ0Z_0\
        );

    \I__7405\ : Odrv4
    port map (
            O => \N__32969\,
            I => \quadWriteZ0Z_0\
        );

    \I__7404\ : InMux
    port map (
            O => \N__32958\,
            I => \N__32955\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__32955\,
            I => \N__32952\
        );

    \I__7402\ : Odrv12
    port map (
            O => \N__32952\,
            I => \MOSIrZ0Z_0\
        );

    \I__7401\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32941\
        );

    \I__7400\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32938\
        );

    \I__7399\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32935\
        );

    \I__7398\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32930\
        );

    \I__7397\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32930\
        );

    \I__7396\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32927\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__32941\,
            I => \N__32923\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__32938\,
            I => \N__32919\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__32935\,
            I => \N__32916\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__32930\,
            I => \N__32911\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__32927\,
            I => \N__32911\
        );

    \I__7390\ : InMux
    port map (
            O => \N__32926\,
            I => \N__32905\
        );

    \I__7389\ : Span4Mux_v
    port map (
            O => \N__32923\,
            I => \N__32902\
        );

    \I__7388\ : InMux
    port map (
            O => \N__32922\,
            I => \N__32899\
        );

    \I__7387\ : Span4Mux_h
    port map (
            O => \N__32919\,
            I => \N__32892\
        );

    \I__7386\ : Span4Mux_h
    port map (
            O => \N__32916\,
            I => \N__32892\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__32911\,
            I => \N__32892\
        );

    \I__7384\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32887\
        );

    \I__7383\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32887\
        );

    \I__7382\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32884\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__32905\,
            I => \data_received_0_repZ0Z2\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__32902\,
            I => \data_received_0_repZ0Z2\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__32899\,
            I => \data_received_0_repZ0Z2\
        );

    \I__7378\ : Odrv4
    port map (
            O => \N__32892\,
            I => \data_received_0_repZ0Z2\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__32887\,
            I => \data_received_0_repZ0Z2\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__32884\,
            I => \data_received_0_repZ0Z2\
        );

    \I__7375\ : InMux
    port map (
            O => \N__32871\,
            I => \N__32868\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__32868\,
            I => \N__32863\
        );

    \I__7373\ : InMux
    port map (
            O => \N__32867\,
            I => \N__32860\
        );

    \I__7372\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32857\
        );

    \I__7371\ : Span4Mux_v
    port map (
            O => \N__32863\,
            I => \N__32854\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__32860\,
            I => \N__32851\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__32857\,
            I => \N__32848\
        );

    \I__7368\ : Odrv4
    port map (
            O => \N__32854\,
            I => \dataRead4_10\
        );

    \I__7367\ : Odrv4
    port map (
            O => \N__32851\,
            I => \dataRead4_10\
        );

    \I__7366\ : Odrv4
    port map (
            O => \N__32848\,
            I => \dataRead4_10\
        );

    \I__7365\ : CascadeMux
    port map (
            O => \N__32841\,
            I => \N__32836\
        );

    \I__7364\ : CascadeMux
    port map (
            O => \N__32840\,
            I => \N__32832\
        );

    \I__7363\ : InMux
    port map (
            O => \N__32839\,
            I => \N__32827\
        );

    \I__7362\ : InMux
    port map (
            O => \N__32836\,
            I => \N__32822\
        );

    \I__7361\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32822\
        );

    \I__7360\ : InMux
    port map (
            O => \N__32832\,
            I => \N__32819\
        );

    \I__7359\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32815\
        );

    \I__7358\ : InMux
    port map (
            O => \N__32830\,
            I => \N__32812\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__32827\,
            I => \N__32807\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__32822\,
            I => \N__32802\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__32819\,
            I => \N__32802\
        );

    \I__7354\ : CascadeMux
    port map (
            O => \N__32818\,
            I => \N__32797\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__32815\,
            I => \N__32794\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__32812\,
            I => \N__32791\
        );

    \I__7351\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32788\
        );

    \I__7350\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32785\
        );

    \I__7349\ : Span4Mux_h
    port map (
            O => \N__32807\,
            I => \N__32780\
        );

    \I__7348\ : Span4Mux_h
    port map (
            O => \N__32802\,
            I => \N__32780\
        );

    \I__7347\ : InMux
    port map (
            O => \N__32801\,
            I => \N__32775\
        );

    \I__7346\ : InMux
    port map (
            O => \N__32800\,
            I => \N__32775\
        );

    \I__7345\ : InMux
    port map (
            O => \N__32797\,
            I => \N__32772\
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__32794\,
            I => \data_received_2_repZ0Z2\
        );

    \I__7343\ : Odrv4
    port map (
            O => \N__32791\,
            I => \data_received_2_repZ0Z2\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__32788\,
            I => \data_received_2_repZ0Z2\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__32785\,
            I => \data_received_2_repZ0Z2\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__32780\,
            I => \data_received_2_repZ0Z2\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__32775\,
            I => \data_received_2_repZ0Z2\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__32772\,
            I => \data_received_2_repZ0Z2\
        );

    \I__7337\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32754\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__32754\,
            I => \QuadInstance0.Quad_RNO_0_0_10\
        );

    \I__7335\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32747\
        );

    \I__7334\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32744\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__32747\,
            I => \QuadInstance0.delayedCh_BZ0Z_1\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__32744\,
            I => \QuadInstance0.delayedCh_BZ0Z_1\
        );

    \I__7331\ : InMux
    port map (
            O => \N__32739\,
            I => \N__32736\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__32736\,
            I => \QuadInstance0.delayedCh_AZ0Z_2\
        );

    \I__7329\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32730\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__32730\,
            I => \N__32726\
        );

    \I__7327\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32723\
        );

    \I__7326\ : Span4Mux_v
    port map (
            O => \N__32726\,
            I => \N__32720\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__32723\,
            I => \N__32717\
        );

    \I__7324\ : Span4Mux_h
    port map (
            O => \N__32720\,
            I => \N__32713\
        );

    \I__7323\ : Span4Mux_v
    port map (
            O => \N__32717\,
            I => \N__32710\
        );

    \I__7322\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32707\
        );

    \I__7321\ : Odrv4
    port map (
            O => \N__32713\,
            I => \dataRead0_1\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__32710\,
            I => \dataRead0_1\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__32707\,
            I => \dataRead0_1\
        );

    \I__7318\ : CascadeMux
    port map (
            O => \N__32700\,
            I => \QuadInstance0.count_enable_cascade_\
        );

    \I__7317\ : CascadeMux
    port map (
            O => \N__32697\,
            I => \N__32694\
        );

    \I__7316\ : InMux
    port map (
            O => \N__32694\,
            I => \N__32691\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__32691\,
            I => \QuadInstance0.Quad_RNIGEBH1Z0Z_1\
        );

    \I__7314\ : CascadeMux
    port map (
            O => \N__32688\,
            I => \N__32684\
        );

    \I__7313\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32680\
        );

    \I__7312\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32675\
        );

    \I__7311\ : InMux
    port map (
            O => \N__32683\,
            I => \N__32675\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__32680\,
            I => \dataRead0_10\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__32675\,
            I => \dataRead0_10\
        );

    \I__7308\ : CascadeMux
    port map (
            O => \N__32670\,
            I => \N__32667\
        );

    \I__7307\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32664\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__32664\,
            I => \QuadInstance0.Quad_RNI0L8Q1Z0Z_10\
        );

    \I__7305\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32658\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__32658\,
            I => \N__32654\
        );

    \I__7303\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32651\
        );

    \I__7302\ : Span4Mux_h
    port map (
            O => \N__32654\,
            I => \N__32645\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__32651\,
            I => \N__32645\
        );

    \I__7300\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32642\
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__32645\,
            I => \dataRead0_2\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__32642\,
            I => \dataRead0_2\
        );

    \I__7297\ : CascadeMux
    port map (
            O => \N__32637\,
            I => \N__32634\
        );

    \I__7296\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32631\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__32631\,
            I => \QuadInstance0.Quad_RNIHFBH1Z0Z_2\
        );

    \I__7294\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32622\
        );

    \I__7293\ : InMux
    port map (
            O => \N__32627\,
            I => \N__32622\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__32622\,
            I => \QuadInstance0.delayedCh_BZ0Z_2\
        );

    \I__7291\ : CascadeMux
    port map (
            O => \N__32619\,
            I => \N__32616\
        );

    \I__7290\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32613\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32610\
        );

    \I__7288\ : Odrv4
    port map (
            O => \N__32610\,
            I => \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_1\
        );

    \I__7287\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32604\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__32604\,
            I => \N__32601\
        );

    \I__7285\ : Odrv4
    port map (
            O => \N__32601\,
            I => \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_1\
        );

    \I__7284\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32595\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__32595\,
            I => \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_1\
        );

    \I__7282\ : CascadeMux
    port map (
            O => \N__32592\,
            I => \N__32563\
        );

    \I__7281\ : CascadeMux
    port map (
            O => \N__32591\,
            I => \N__32560\
        );

    \I__7280\ : CascadeMux
    port map (
            O => \N__32590\,
            I => \N__32557\
        );

    \I__7279\ : CascadeMux
    port map (
            O => \N__32589\,
            I => \N__32554\
        );

    \I__7278\ : CascadeMux
    port map (
            O => \N__32588\,
            I => \N__32551\
        );

    \I__7277\ : CascadeMux
    port map (
            O => \N__32587\,
            I => \N__32548\
        );

    \I__7276\ : CascadeMux
    port map (
            O => \N__32586\,
            I => \N__32545\
        );

    \I__7275\ : CascadeMux
    port map (
            O => \N__32585\,
            I => \N__32535\
        );

    \I__7274\ : CascadeMux
    port map (
            O => \N__32584\,
            I => \N__32531\
        );

    \I__7273\ : CascadeMux
    port map (
            O => \N__32583\,
            I => \N__32528\
        );

    \I__7272\ : CascadeMux
    port map (
            O => \N__32582\,
            I => \N__32525\
        );

    \I__7271\ : CascadeMux
    port map (
            O => \N__32581\,
            I => \N__32522\
        );

    \I__7270\ : CascadeMux
    port map (
            O => \N__32580\,
            I => \N__32519\
        );

    \I__7269\ : CascadeMux
    port map (
            O => \N__32579\,
            I => \N__32515\
        );

    \I__7268\ : CascadeMux
    port map (
            O => \N__32578\,
            I => \N__32512\
        );

    \I__7267\ : CascadeMux
    port map (
            O => \N__32577\,
            I => \N__32509\
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__32576\,
            I => \N__32506\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__32575\,
            I => \N__32503\
        );

    \I__7264\ : CascadeMux
    port map (
            O => \N__32574\,
            I => \N__32500\
        );

    \I__7263\ : CascadeMux
    port map (
            O => \N__32573\,
            I => \N__32497\
        );

    \I__7262\ : CascadeMux
    port map (
            O => \N__32572\,
            I => \N__32491\
        );

    \I__7261\ : CascadeMux
    port map (
            O => \N__32571\,
            I => \N__32488\
        );

    \I__7260\ : CascadeMux
    port map (
            O => \N__32570\,
            I => \N__32485\
        );

    \I__7259\ : CascadeMux
    port map (
            O => \N__32569\,
            I => \N__32482\
        );

    \I__7258\ : CascadeMux
    port map (
            O => \N__32568\,
            I => \N__32479\
        );

    \I__7257\ : CascadeMux
    port map (
            O => \N__32567\,
            I => \N__32476\
        );

    \I__7256\ : CascadeMux
    port map (
            O => \N__32566\,
            I => \N__32473\
        );

    \I__7255\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32457\
        );

    \I__7254\ : InMux
    port map (
            O => \N__32560\,
            I => \N__32457\
        );

    \I__7253\ : InMux
    port map (
            O => \N__32557\,
            I => \N__32457\
        );

    \I__7252\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32457\
        );

    \I__7251\ : InMux
    port map (
            O => \N__32551\,
            I => \N__32450\
        );

    \I__7250\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32450\
        );

    \I__7249\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32450\
        );

    \I__7248\ : CascadeMux
    port map (
            O => \N__32544\,
            I => \N__32447\
        );

    \I__7247\ : CascadeMux
    port map (
            O => \N__32543\,
            I => \N__32444\
        );

    \I__7246\ : CascadeMux
    port map (
            O => \N__32542\,
            I => \N__32441\
        );

    \I__7245\ : CascadeMux
    port map (
            O => \N__32541\,
            I => \N__32438\
        );

    \I__7244\ : CascadeMux
    port map (
            O => \N__32540\,
            I => \N__32435\
        );

    \I__7243\ : CascadeMux
    port map (
            O => \N__32539\,
            I => \N__32432\
        );

    \I__7242\ : CascadeMux
    port map (
            O => \N__32538\,
            I => \N__32429\
        );

    \I__7241\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32418\
        );

    \I__7240\ : InMux
    port map (
            O => \N__32534\,
            I => \N__32418\
        );

    \I__7239\ : InMux
    port map (
            O => \N__32531\,
            I => \N__32418\
        );

    \I__7238\ : InMux
    port map (
            O => \N__32528\,
            I => \N__32418\
        );

    \I__7237\ : InMux
    port map (
            O => \N__32525\,
            I => \N__32418\
        );

    \I__7236\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32413\
        );

    \I__7235\ : InMux
    port map (
            O => \N__32519\,
            I => \N__32413\
        );

    \I__7234\ : CascadeMux
    port map (
            O => \N__32518\,
            I => \N__32407\
        );

    \I__7233\ : InMux
    port map (
            O => \N__32515\,
            I => \N__32398\
        );

    \I__7232\ : InMux
    port map (
            O => \N__32512\,
            I => \N__32398\
        );

    \I__7231\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32398\
        );

    \I__7230\ : InMux
    port map (
            O => \N__32506\,
            I => \N__32398\
        );

    \I__7229\ : InMux
    port map (
            O => \N__32503\,
            I => \N__32391\
        );

    \I__7228\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32391\
        );

    \I__7227\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32391\
        );

    \I__7226\ : CascadeMux
    port map (
            O => \N__32496\,
            I => \N__32387\
        );

    \I__7225\ : CascadeMux
    port map (
            O => \N__32495\,
            I => \N__32384\
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__32494\,
            I => \N__32379\
        );

    \I__7223\ : InMux
    port map (
            O => \N__32491\,
            I => \N__32370\
        );

    \I__7222\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32370\
        );

    \I__7221\ : InMux
    port map (
            O => \N__32485\,
            I => \N__32370\
        );

    \I__7220\ : InMux
    port map (
            O => \N__32482\,
            I => \N__32370\
        );

    \I__7219\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32363\
        );

    \I__7218\ : InMux
    port map (
            O => \N__32476\,
            I => \N__32363\
        );

    \I__7217\ : InMux
    port map (
            O => \N__32473\,
            I => \N__32363\
        );

    \I__7216\ : CascadeMux
    port map (
            O => \N__32472\,
            I => \N__32360\
        );

    \I__7215\ : CascadeMux
    port map (
            O => \N__32471\,
            I => \N__32357\
        );

    \I__7214\ : CascadeMux
    port map (
            O => \N__32470\,
            I => \N__32354\
        );

    \I__7213\ : CascadeMux
    port map (
            O => \N__32469\,
            I => \N__32351\
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__32468\,
            I => \N__32348\
        );

    \I__7211\ : CascadeMux
    port map (
            O => \N__32467\,
            I => \N__32345\
        );

    \I__7210\ : CascadeMux
    port map (
            O => \N__32466\,
            I => \N__32342\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__32457\,
            I => \N__32339\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__32450\,
            I => \N__32336\
        );

    \I__7207\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32327\
        );

    \I__7206\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32327\
        );

    \I__7205\ : InMux
    port map (
            O => \N__32441\,
            I => \N__32327\
        );

    \I__7204\ : InMux
    port map (
            O => \N__32438\,
            I => \N__32327\
        );

    \I__7203\ : InMux
    port map (
            O => \N__32435\,
            I => \N__32320\
        );

    \I__7202\ : InMux
    port map (
            O => \N__32432\,
            I => \N__32320\
        );

    \I__7201\ : InMux
    port map (
            O => \N__32429\,
            I => \N__32320\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32315\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__32413\,
            I => \N__32315\
        );

    \I__7198\ : CascadeMux
    port map (
            O => \N__32412\,
            I => \N__32311\
        );

    \I__7197\ : CascadeMux
    port map (
            O => \N__32411\,
            I => \N__32308\
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__32410\,
            I => \N__32302\
        );

    \I__7195\ : InMux
    port map (
            O => \N__32407\,
            I => \N__32299\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__32398\,
            I => \N__32294\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__32391\,
            I => \N__32294\
        );

    \I__7192\ : InMux
    port map (
            O => \N__32390\,
            I => \N__32281\
        );

    \I__7191\ : InMux
    port map (
            O => \N__32387\,
            I => \N__32281\
        );

    \I__7190\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32281\
        );

    \I__7189\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32281\
        );

    \I__7188\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32281\
        );

    \I__7187\ : InMux
    port map (
            O => \N__32379\,
            I => \N__32281\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__32370\,
            I => \N__32276\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__32363\,
            I => \N__32276\
        );

    \I__7184\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32267\
        );

    \I__7183\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32267\
        );

    \I__7182\ : InMux
    port map (
            O => \N__32354\,
            I => \N__32267\
        );

    \I__7181\ : InMux
    port map (
            O => \N__32351\,
            I => \N__32267\
        );

    \I__7180\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32260\
        );

    \I__7179\ : InMux
    port map (
            O => \N__32345\,
            I => \N__32260\
        );

    \I__7178\ : InMux
    port map (
            O => \N__32342\,
            I => \N__32260\
        );

    \I__7177\ : Span4Mux_v
    port map (
            O => \N__32339\,
            I => \N__32255\
        );

    \I__7176\ : Span4Mux_v
    port map (
            O => \N__32336\,
            I => \N__32255\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__32327\,
            I => \N__32250\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__32320\,
            I => \N__32250\
        );

    \I__7173\ : Span4Mux_v
    port map (
            O => \N__32315\,
            I => \N__32247\
        );

    \I__7172\ : InMux
    port map (
            O => \N__32314\,
            I => \N__32232\
        );

    \I__7171\ : InMux
    port map (
            O => \N__32311\,
            I => \N__32232\
        );

    \I__7170\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32232\
        );

    \I__7169\ : InMux
    port map (
            O => \N__32307\,
            I => \N__32232\
        );

    \I__7168\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32232\
        );

    \I__7167\ : InMux
    port map (
            O => \N__32305\,
            I => \N__32232\
        );

    \I__7166\ : InMux
    port map (
            O => \N__32302\,
            I => \N__32232\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__32299\,
            I => \N__32229\
        );

    \I__7164\ : Span4Mux_h
    port map (
            O => \N__32294\,
            I => \N__32224\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__32281\,
            I => \N__32224\
        );

    \I__7162\ : Span4Mux_h
    port map (
            O => \N__32276\,
            I => \N__32221\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__32267\,
            I => \N__32216\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__32260\,
            I => \N__32216\
        );

    \I__7159\ : Span4Mux_h
    port map (
            O => \N__32255\,
            I => \N__32211\
        );

    \I__7158\ : Span4Mux_h
    port map (
            O => \N__32250\,
            I => \N__32211\
        );

    \I__7157\ : Sp12to4
    port map (
            O => \N__32247\,
            I => \N__32208\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__32232\,
            I => \N__32205\
        );

    \I__7155\ : Span4Mux_v
    port map (
            O => \N__32229\,
            I => \N__32202\
        );

    \I__7154\ : Span4Mux_v
    port map (
            O => \N__32224\,
            I => \N__32199\
        );

    \I__7153\ : Span4Mux_v
    port map (
            O => \N__32221\,
            I => \N__32194\
        );

    \I__7152\ : Span4Mux_h
    port map (
            O => \N__32216\,
            I => \N__32194\
        );

    \I__7151\ : Span4Mux_v
    port map (
            O => \N__32211\,
            I => \N__32191\
        );

    \I__7150\ : Span12Mux_h
    port map (
            O => \N__32208\,
            I => \N__32186\
        );

    \I__7149\ : Sp12to4
    port map (
            O => \N__32205\,
            I => \N__32186\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__32202\,
            I => \N__32179\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__32199\,
            I => \N__32179\
        );

    \I__7146\ : Span4Mux_h
    port map (
            O => \N__32194\,
            I => \N__32179\
        );

    \I__7145\ : Odrv4
    port map (
            O => \N__32191\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7144\ : Odrv12
    port map (
            O => \N__32186\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__32179\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7142\ : CascadeMux
    port map (
            O => \N__32172\,
            I => \N__32169\
        );

    \I__7141\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32166\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__32166\,
            I => \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_1\
        );

    \I__7139\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32160\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__32160\,
            I => \N__32157\
        );

    \I__7137\ : Odrv12
    port map (
            O => \N__32157\,
            I => \PWMInstance2.un1_periodCounter12_1_0_a2_0\
        );

    \I__7136\ : InMux
    port map (
            O => \N__32154\,
            I => \bfn_17_15_0_\
        );

    \I__7135\ : IoInMux
    port map (
            O => \N__32151\,
            I => \N__32148\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__32148\,
            I => \N__32145\
        );

    \I__7133\ : Span4Mux_s1_v
    port map (
            O => \N__32145\,
            I => \N__32142\
        );

    \I__7132\ : Span4Mux_v
    port map (
            O => \N__32142\,
            I => \N__32138\
        );

    \I__7131\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32135\
        );

    \I__7130\ : Odrv4
    port map (
            O => \N__32138\,
            I => \PWM2_c\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__32135\,
            I => \PWM2_c\
        );

    \I__7128\ : InMux
    port map (
            O => \N__32130\,
            I => \N__32127\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__32127\,
            I => \MOSI_c\
        );

    \I__7126\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32121\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__32121\,
            I => \ch1_A_c\
        );

    \I__7124\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32115\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__32115\,
            I => \N__32112\
        );

    \I__7122\ : Span4Mux_h
    port map (
            O => \N__32112\,
            I => \N__32109\
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__32109\,
            I => \QuadInstance1.delayedCh_AZ0Z_0\
        );

    \I__7120\ : InMux
    port map (
            O => \N__32106\,
            I => \N__32103\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32100\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__32100\,
            I => \N__32097\
        );

    \I__7117\ : Span4Mux_h
    port map (
            O => \N__32097\,
            I => \N__32094\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__32094\,
            I => \QuadInstance0.delayedCh_AZ0Z_0\
        );

    \I__7115\ : InMux
    port map (
            O => \N__32091\,
            I => \N__32088\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__32088\,
            I => \N__32079\
        );

    \I__7113\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32074\
        );

    \I__7112\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32074\
        );

    \I__7111\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32069\
        );

    \I__7110\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32066\
        );

    \I__7109\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32063\
        );

    \I__7108\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32060\
        );

    \I__7107\ : Span4Mux_v
    port map (
            O => \N__32079\,
            I => \N__32057\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__32074\,
            I => \N__32054\
        );

    \I__7105\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32051\
        );

    \I__7104\ : InMux
    port map (
            O => \N__32072\,
            I => \N__32047\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__32069\,
            I => \N__32044\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__32066\,
            I => \N__32040\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__32063\,
            I => \N__32037\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__32060\,
            I => \N__32034\
        );

    \I__7099\ : Span4Mux_h
    port map (
            O => \N__32057\,
            I => \N__32026\
        );

    \I__7098\ : Span4Mux_v
    port map (
            O => \N__32054\,
            I => \N__32026\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__32051\,
            I => \N__32026\
        );

    \I__7096\ : InMux
    port map (
            O => \N__32050\,
            I => \N__32023\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__32047\,
            I => \N__32017\
        );

    \I__7094\ : Span4Mux_h
    port map (
            O => \N__32044\,
            I => \N__32014\
        );

    \I__7093\ : InMux
    port map (
            O => \N__32043\,
            I => \N__32011\
        );

    \I__7092\ : Span4Mux_h
    port map (
            O => \N__32040\,
            I => \N__32008\
        );

    \I__7091\ : Span4Mux_h
    port map (
            O => \N__32037\,
            I => \N__32005\
        );

    \I__7090\ : Span4Mux_v
    port map (
            O => \N__32034\,
            I => \N__32002\
        );

    \I__7089\ : InMux
    port map (
            O => \N__32033\,
            I => \N__31999\
        );

    \I__7088\ : Span4Mux_h
    port map (
            O => \N__32026\,
            I => \N__31994\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__32023\,
            I => \N__31994\
        );

    \I__7086\ : InMux
    port map (
            O => \N__32022\,
            I => \N__31989\
        );

    \I__7085\ : InMux
    port map (
            O => \N__32021\,
            I => \N__31989\
        );

    \I__7084\ : InMux
    port map (
            O => \N__32020\,
            I => \N__31986\
        );

    \I__7083\ : Span4Mux_h
    port map (
            O => \N__32017\,
            I => \N__31978\
        );

    \I__7082\ : Span4Mux_h
    port map (
            O => \N__32014\,
            I => \N__31978\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__32011\,
            I => \N__31978\
        );

    \I__7080\ : Span4Mux_h
    port map (
            O => \N__32008\,
            I => \N__31973\
        );

    \I__7079\ : Span4Mux_v
    port map (
            O => \N__32005\,
            I => \N__31973\
        );

    \I__7078\ : Span4Mux_h
    port map (
            O => \N__32002\,
            I => \N__31970\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__31999\,
            I => \N__31967\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__31994\,
            I => \N__31964\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__31989\,
            I => \N__31959\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__31986\,
            I => \N__31959\
        );

    \I__7073\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31956\
        );

    \I__7072\ : Span4Mux_v
    port map (
            O => \N__31978\,
            I => \N__31951\
        );

    \I__7071\ : Span4Mux_h
    port map (
            O => \N__31973\,
            I => \N__31951\
        );

    \I__7070\ : Span4Mux_h
    port map (
            O => \N__31970\,
            I => \N__31942\
        );

    \I__7069\ : Span4Mux_h
    port map (
            O => \N__31967\,
            I => \N__31942\
        );

    \I__7068\ : Span4Mux_h
    port map (
            O => \N__31964\,
            I => \N__31942\
        );

    \I__7067\ : Span4Mux_h
    port map (
            O => \N__31959\,
            I => \N__31942\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__31956\,
            I => \dataWriteZ0Z_3\
        );

    \I__7065\ : Odrv4
    port map (
            O => \N__31951\,
            I => \dataWriteZ0Z_3\
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__31942\,
            I => \dataWriteZ0Z_3\
        );

    \I__7063\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31932\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__31932\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_3\
        );

    \I__7061\ : InMux
    port map (
            O => \N__31929\,
            I => \N__31926\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__31926\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_14\
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__31923\,
            I => \N__31920\
        );

    \I__7058\ : InMux
    port map (
            O => \N__31920\,
            I => \N__31913\
        );

    \I__7057\ : CascadeMux
    port map (
            O => \N__31919\,
            I => \N__31910\
        );

    \I__7056\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31905\
        );

    \I__7055\ : CascadeMux
    port map (
            O => \N__31917\,
            I => \N__31900\
        );

    \I__7054\ : CascadeMux
    port map (
            O => \N__31916\,
            I => \N__31897\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__31913\,
            I => \N__31891\
        );

    \I__7052\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31888\
        );

    \I__7051\ : CascadeMux
    port map (
            O => \N__31909\,
            I => \N__31885\
        );

    \I__7050\ : CascadeMux
    port map (
            O => \N__31908\,
            I => \N__31882\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__31905\,
            I => \N__31879\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31904\,
            I => \N__31875\
        );

    \I__7047\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31872\
        );

    \I__7046\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31868\
        );

    \I__7045\ : InMux
    port map (
            O => \N__31897\,
            I => \N__31865\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__31896\,
            I => \N__31862\
        );

    \I__7043\ : CascadeMux
    port map (
            O => \N__31895\,
            I => \N__31859\
        );

    \I__7042\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31854\
        );

    \I__7041\ : Span4Mux_h
    port map (
            O => \N__31891\,
            I => \N__31849\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__31888\,
            I => \N__31849\
        );

    \I__7039\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31846\
        );

    \I__7038\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31843\
        );

    \I__7037\ : Span4Mux_v
    port map (
            O => \N__31879\,
            I => \N__31840\
        );

    \I__7036\ : InMux
    port map (
            O => \N__31878\,
            I => \N__31837\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__31875\,
            I => \N__31832\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__31872\,
            I => \N__31832\
        );

    \I__7033\ : InMux
    port map (
            O => \N__31871\,
            I => \N__31829\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__31868\,
            I => \N__31826\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__31865\,
            I => \N__31823\
        );

    \I__7030\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31820\
        );

    \I__7029\ : InMux
    port map (
            O => \N__31859\,
            I => \N__31817\
        );

    \I__7028\ : InMux
    port map (
            O => \N__31858\,
            I => \N__31814\
        );

    \I__7027\ : InMux
    port map (
            O => \N__31857\,
            I => \N__31811\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__31854\,
            I => \N__31808\
        );

    \I__7025\ : Span4Mux_v
    port map (
            O => \N__31849\,
            I => \N__31801\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__31846\,
            I => \N__31801\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__31843\,
            I => \N__31801\
        );

    \I__7022\ : Span4Mux_h
    port map (
            O => \N__31840\,
            I => \N__31798\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__31837\,
            I => \N__31795\
        );

    \I__7020\ : Span4Mux_v
    port map (
            O => \N__31832\,
            I => \N__31792\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__31829\,
            I => \N__31789\
        );

    \I__7018\ : Span4Mux_v
    port map (
            O => \N__31826\,
            I => \N__31786\
        );

    \I__7017\ : Span4Mux_h
    port map (
            O => \N__31823\,
            I => \N__31779\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__31820\,
            I => \N__31779\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__31817\,
            I => \N__31779\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__31814\,
            I => \N__31776\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__31811\,
            I => \N__31773\
        );

    \I__7012\ : Span4Mux_v
    port map (
            O => \N__31808\,
            I => \N__31768\
        );

    \I__7011\ : Span4Mux_v
    port map (
            O => \N__31801\,
            I => \N__31768\
        );

    \I__7010\ : Span4Mux_v
    port map (
            O => \N__31798\,
            I => \N__31765\
        );

    \I__7009\ : Span4Mux_v
    port map (
            O => \N__31795\,
            I => \N__31758\
        );

    \I__7008\ : Span4Mux_h
    port map (
            O => \N__31792\,
            I => \N__31758\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__31789\,
            I => \N__31758\
        );

    \I__7006\ : Span4Mux_h
    port map (
            O => \N__31786\,
            I => \N__31753\
        );

    \I__7005\ : Span4Mux_v
    port map (
            O => \N__31779\,
            I => \N__31753\
        );

    \I__7004\ : Span4Mux_v
    port map (
            O => \N__31776\,
            I => \N__31746\
        );

    \I__7003\ : Span4Mux_v
    port map (
            O => \N__31773\,
            I => \N__31746\
        );

    \I__7002\ : Span4Mux_h
    port map (
            O => \N__31768\,
            I => \N__31746\
        );

    \I__7001\ : Odrv4
    port map (
            O => \N__31765\,
            I => \dataWriteZ0Z_15\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__31758\,
            I => \dataWriteZ0Z_15\
        );

    \I__6999\ : Odrv4
    port map (
            O => \N__31753\,
            I => \dataWriteZ0Z_15\
        );

    \I__6998\ : Odrv4
    port map (
            O => \N__31746\,
            I => \dataWriteZ0Z_15\
        );

    \I__6997\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31734\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__31734\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_15\
        );

    \I__6995\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31728\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__31725\,
            I => \N__31722\
        );

    \I__6992\ : Odrv4
    port map (
            O => \N__31722\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_13\
        );

    \I__6991\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31716\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__31716\,
            I => \N__31713\
        );

    \I__6989\ : Odrv4
    port map (
            O => \N__31713\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_12\
        );

    \I__6988\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__31707\,
            I => \N__31704\
        );

    \I__6986\ : Odrv12
    port map (
            O => \N__31704\,
            I => \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_1\
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__31701\,
            I => \N__31698\
        );

    \I__6984\ : InMux
    port map (
            O => \N__31698\,
            I => \N__31695\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__31695\,
            I => \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_1\
        );

    \I__6982\ : InMux
    port map (
            O => \N__31692\,
            I => \N__31683\
        );

    \I__6981\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31683\
        );

    \I__6980\ : InMux
    port map (
            O => \N__31690\,
            I => \N__31683\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__31683\,
            I => \N__31680\
        );

    \I__6978\ : Odrv4
    port map (
            O => \N__31680\,
            I => \pwmWriteZ0Z_2\
        );

    \I__6977\ : InMux
    port map (
            O => \N__31677\,
            I => \N__31671\
        );

    \I__6976\ : InMux
    port map (
            O => \N__31676\,
            I => \N__31671\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__31671\,
            I => \N__31668\
        );

    \I__6974\ : Odrv12
    port map (
            O => \N__31668\,
            I => \pwmWrite_fastZ0Z_2\
        );

    \I__6973\ : CascadeMux
    port map (
            O => \N__31665\,
            I => \N__31661\
        );

    \I__6972\ : CascadeMux
    port map (
            O => \N__31664\,
            I => \N__31658\
        );

    \I__6971\ : InMux
    port map (
            O => \N__31661\,
            I => \N__31647\
        );

    \I__6970\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31647\
        );

    \I__6969\ : InMux
    port map (
            O => \N__31657\,
            I => \N__31647\
        );

    \I__6968\ : InMux
    port map (
            O => \N__31656\,
            I => \N__31647\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__31647\,
            I => \PWMInstance2.clkCountZ0Z_1\
        );

    \I__6966\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31632\
        );

    \I__6965\ : InMux
    port map (
            O => \N__31643\,
            I => \N__31632\
        );

    \I__6964\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31632\
        );

    \I__6963\ : InMux
    port map (
            O => \N__31641\,
            I => \N__31632\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__31632\,
            I => \PWMInstance2.clkCountZ0Z_0\
        );

    \I__6961\ : CascadeMux
    port map (
            O => \N__31629\,
            I => \PWMInstance2.un1_periodCounter12_1_0_a2_0_6_cascade_\
        );

    \I__6960\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31623\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__31623\,
            I => \PWMInstance2.un1_periodCounter12_1_0_a2_0_9\
        );

    \I__6958\ : CascadeMux
    port map (
            O => \N__31620\,
            I => \PWMInstance2.un1_periodCounter12_1_0_a2_0_14_cascade_\
        );

    \I__6957\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31614\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__31614\,
            I => \N__31611\
        );

    \I__6955\ : Odrv4
    port map (
            O => \N__31611\,
            I => \PWMInstance2.un1_periodCounter12_1_0_a2_0_10\
        );

    \I__6954\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31605\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__31605\,
            I => \N__31600\
        );

    \I__6952\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31597\
        );

    \I__6951\ : InMux
    port map (
            O => \N__31603\,
            I => \N__31594\
        );

    \I__6950\ : Span4Mux_s2_v
    port map (
            O => \N__31600\,
            I => \N__31580\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__31597\,
            I => \N__31577\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__31594\,
            I => \N__31574\
        );

    \I__6947\ : InMux
    port map (
            O => \N__31593\,
            I => \N__31571\
        );

    \I__6946\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31568\
        );

    \I__6945\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31565\
        );

    \I__6944\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31560\
        );

    \I__6943\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31560\
        );

    \I__6942\ : InMux
    port map (
            O => \N__31588\,
            I => \N__31555\
        );

    \I__6941\ : InMux
    port map (
            O => \N__31587\,
            I => \N__31555\
        );

    \I__6940\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31550\
        );

    \I__6939\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31550\
        );

    \I__6938\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31547\
        );

    \I__6937\ : InMux
    port map (
            O => \N__31583\,
            I => \N__31544\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__31580\,
            I => \N__31539\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__31577\,
            I => \N__31534\
        );

    \I__6934\ : Span4Mux_v
    port map (
            O => \N__31574\,
            I => \N__31534\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__31571\,
            I => \N__31531\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31528\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__31565\,
            I => \N__31525\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__31560\,
            I => \N__31520\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__31555\,
            I => \N__31520\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__31550\,
            I => \N__31517\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__31547\,
            I => \N__31512\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__31544\,
            I => \N__31512\
        );

    \I__6925\ : InMux
    port map (
            O => \N__31543\,
            I => \N__31509\
        );

    \I__6924\ : InMux
    port map (
            O => \N__31542\,
            I => \N__31506\
        );

    \I__6923\ : Span4Mux_v
    port map (
            O => \N__31539\,
            I => \N__31501\
        );

    \I__6922\ : Span4Mux_h
    port map (
            O => \N__31534\,
            I => \N__31501\
        );

    \I__6921\ : Span4Mux_h
    port map (
            O => \N__31531\,
            I => \N__31498\
        );

    \I__6920\ : Span4Mux_v
    port map (
            O => \N__31528\,
            I => \N__31493\
        );

    \I__6919\ : Span4Mux_h
    port map (
            O => \N__31525\,
            I => \N__31493\
        );

    \I__6918\ : Span4Mux_h
    port map (
            O => \N__31520\,
            I => \N__31488\
        );

    \I__6917\ : Span4Mux_h
    port map (
            O => \N__31517\,
            I => \N__31488\
        );

    \I__6916\ : Span4Mux_h
    port map (
            O => \N__31512\,
            I => \N__31483\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__31509\,
            I => \N__31483\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__31506\,
            I => \N__31480\
        );

    \I__6913\ : Span4Mux_h
    port map (
            O => \N__31501\,
            I => \N__31477\
        );

    \I__6912\ : Span4Mux_h
    port map (
            O => \N__31498\,
            I => \N__31474\
        );

    \I__6911\ : Span4Mux_h
    port map (
            O => \N__31493\,
            I => \N__31469\
        );

    \I__6910\ : Span4Mux_v
    port map (
            O => \N__31488\,
            I => \N__31469\
        );

    \I__6909\ : Span4Mux_v
    port map (
            O => \N__31483\,
            I => \N__31464\
        );

    \I__6908\ : Span4Mux_h
    port map (
            O => \N__31480\,
            I => \N__31464\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__31477\,
            I => \dataWriteZ0Z_2\
        );

    \I__6906\ : Odrv4
    port map (
            O => \N__31474\,
            I => \dataWriteZ0Z_2\
        );

    \I__6905\ : Odrv4
    port map (
            O => \N__31469\,
            I => \dataWriteZ0Z_2\
        );

    \I__6904\ : Odrv4
    port map (
            O => \N__31464\,
            I => \dataWriteZ0Z_2\
        );

    \I__6903\ : CascadeMux
    port map (
            O => \N__31455\,
            I => \N__31452\
        );

    \I__6902\ : InMux
    port map (
            O => \N__31452\,
            I => \N__31449\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__31449\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_2\
        );

    \I__6900\ : InMux
    port map (
            O => \N__31446\,
            I => \N__31443\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__31443\,
            I => \OutReg_0_sqmuxa_0_a2_3_a2_2\
        );

    \I__6898\ : CascadeMux
    port map (
            O => \N__31440\,
            I => \N__31431\
        );

    \I__6897\ : CascadeMux
    port map (
            O => \N__31439\,
            I => \N__31426\
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__31438\,
            I => \N__31423\
        );

    \I__6895\ : InMux
    port map (
            O => \N__31437\,
            I => \N__31419\
        );

    \I__6894\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31416\
        );

    \I__6893\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31413\
        );

    \I__6892\ : CascadeMux
    port map (
            O => \N__31434\,
            I => \N__31408\
        );

    \I__6891\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31404\
        );

    \I__6890\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31395\
        );

    \I__6889\ : InMux
    port map (
            O => \N__31429\,
            I => \N__31395\
        );

    \I__6888\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31395\
        );

    \I__6887\ : InMux
    port map (
            O => \N__31423\,
            I => \N__31395\
        );

    \I__6886\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31392\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__31419\,
            I => \N__31389\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__31416\,
            I => \N__31386\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__31413\,
            I => \N__31383\
        );

    \I__6882\ : InMux
    port map (
            O => \N__31412\,
            I => \N__31379\
        );

    \I__6881\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31375\
        );

    \I__6880\ : InMux
    port map (
            O => \N__31408\,
            I => \N__31369\
        );

    \I__6879\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31369\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__31404\,
            I => \N__31364\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__31395\,
            I => \N__31364\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__31392\,
            I => \N__31361\
        );

    \I__6875\ : Span4Mux_v
    port map (
            O => \N__31389\,
            I => \N__31358\
        );

    \I__6874\ : Span4Mux_v
    port map (
            O => \N__31386\,
            I => \N__31355\
        );

    \I__6873\ : Span4Mux_v
    port map (
            O => \N__31383\,
            I => \N__31352\
        );

    \I__6872\ : InMux
    port map (
            O => \N__31382\,
            I => \N__31349\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__31379\,
            I => \N__31346\
        );

    \I__6870\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31343\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__31375\,
            I => \N__31340\
        );

    \I__6868\ : InMux
    port map (
            O => \N__31374\,
            I => \N__31337\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__31369\,
            I => \N__31332\
        );

    \I__6866\ : Span4Mux_h
    port map (
            O => \N__31364\,
            I => \N__31332\
        );

    \I__6865\ : Span4Mux_v
    port map (
            O => \N__31361\,
            I => \N__31325\
        );

    \I__6864\ : Span4Mux_h
    port map (
            O => \N__31358\,
            I => \N__31325\
        );

    \I__6863\ : Span4Mux_h
    port map (
            O => \N__31355\,
            I => \N__31325\
        );

    \I__6862\ : Span4Mux_v
    port map (
            O => \N__31352\,
            I => \N__31322\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__31349\,
            I => \N__31317\
        );

    \I__6860\ : Span4Mux_v
    port map (
            O => \N__31346\,
            I => \N__31317\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__31343\,
            I => \N__31314\
        );

    \I__6858\ : Span4Mux_h
    port map (
            O => \N__31340\,
            I => \N__31311\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__31337\,
            I => \N__31308\
        );

    \I__6856\ : Span4Mux_v
    port map (
            O => \N__31332\,
            I => \N__31303\
        );

    \I__6855\ : Span4Mux_h
    port map (
            O => \N__31325\,
            I => \N__31303\
        );

    \I__6854\ : Span4Mux_h
    port map (
            O => \N__31322\,
            I => \N__31298\
        );

    \I__6853\ : Span4Mux_h
    port map (
            O => \N__31317\,
            I => \N__31298\
        );

    \I__6852\ : Odrv12
    port map (
            O => \N__31314\,
            I => \dataWriteZ0Z_0\
        );

    \I__6851\ : Odrv4
    port map (
            O => \N__31311\,
            I => \dataWriteZ0Z_0\
        );

    \I__6850\ : Odrv12
    port map (
            O => \N__31308\,
            I => \dataWriteZ0Z_0\
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__31303\,
            I => \dataWriteZ0Z_0\
        );

    \I__6848\ : Odrv4
    port map (
            O => \N__31298\,
            I => \dataWriteZ0Z_0\
        );

    \I__6847\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31284\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__31284\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_0\
        );

    \I__6845\ : InMux
    port map (
            O => \N__31281\,
            I => \N__31275\
        );

    \I__6844\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31272\
        );

    \I__6843\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31268\
        );

    \I__6842\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31265\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__31275\,
            I => \N__31261\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__31272\,
            I => \N__31258\
        );

    \I__6839\ : InMux
    port map (
            O => \N__31271\,
            I => \N__31253\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__31268\,
            I => \N__31249\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__31265\,
            I => \N__31244\
        );

    \I__6836\ : InMux
    port map (
            O => \N__31264\,
            I => \N__31241\
        );

    \I__6835\ : Span4Mux_v
    port map (
            O => \N__31261\,
            I => \N__31236\
        );

    \I__6834\ : Span4Mux_v
    port map (
            O => \N__31258\,
            I => \N__31233\
        );

    \I__6833\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31230\
        );

    \I__6832\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31227\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__31253\,
            I => \N__31224\
        );

    \I__6830\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31221\
        );

    \I__6829\ : Span4Mux_h
    port map (
            O => \N__31249\,
            I => \N__31215\
        );

    \I__6828\ : InMux
    port map (
            O => \N__31248\,
            I => \N__31212\
        );

    \I__6827\ : InMux
    port map (
            O => \N__31247\,
            I => \N__31209\
        );

    \I__6826\ : Span4Mux_v
    port map (
            O => \N__31244\,
            I => \N__31206\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__31241\,
            I => \N__31203\
        );

    \I__6824\ : InMux
    port map (
            O => \N__31240\,
            I => \N__31200\
        );

    \I__6823\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31197\
        );

    \I__6822\ : Span4Mux_h
    port map (
            O => \N__31236\,
            I => \N__31190\
        );

    \I__6821\ : Span4Mux_h
    port map (
            O => \N__31233\,
            I => \N__31190\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__31230\,
            I => \N__31190\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31187\
        );

    \I__6818\ : Span4Mux_s2_v
    port map (
            O => \N__31224\,
            I => \N__31182\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__31221\,
            I => \N__31182\
        );

    \I__6816\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31175\
        );

    \I__6815\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31175\
        );

    \I__6814\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31175\
        );

    \I__6813\ : Span4Mux_v
    port map (
            O => \N__31215\,
            I => \N__31168\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__31212\,
            I => \N__31168\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__31209\,
            I => \N__31168\
        );

    \I__6810\ : Span4Mux_h
    port map (
            O => \N__31206\,
            I => \N__31163\
        );

    \I__6809\ : Span4Mux_v
    port map (
            O => \N__31203\,
            I => \N__31163\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31158\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__31197\,
            I => \N__31158\
        );

    \I__6806\ : Span4Mux_v
    port map (
            O => \N__31190\,
            I => \N__31153\
        );

    \I__6805\ : Span4Mux_h
    port map (
            O => \N__31187\,
            I => \N__31153\
        );

    \I__6804\ : Span4Mux_v
    port map (
            O => \N__31182\,
            I => \N__31146\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__31175\,
            I => \N__31146\
        );

    \I__6802\ : Span4Mux_h
    port map (
            O => \N__31168\,
            I => \N__31146\
        );

    \I__6801\ : Odrv4
    port map (
            O => \N__31163\,
            I => \dataWriteZ0Z_1\
        );

    \I__6800\ : Odrv12
    port map (
            O => \N__31158\,
            I => \dataWriteZ0Z_1\
        );

    \I__6799\ : Odrv4
    port map (
            O => \N__31153\,
            I => \dataWriteZ0Z_1\
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__31146\,
            I => \dataWriteZ0Z_1\
        );

    \I__6797\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__31134\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_1\
        );

    \I__6795\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31128\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__31128\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_7\
        );

    \I__6793\ : InMux
    port map (
            O => \N__31125\,
            I => \N__31121\
        );

    \I__6792\ : InMux
    port map (
            O => \N__31124\,
            I => \N__31115\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__31121\,
            I => \N__31104\
        );

    \I__6790\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31101\
        );

    \I__6789\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31098\
        );

    \I__6788\ : InMux
    port map (
            O => \N__31118\,
            I => \N__31095\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__31115\,
            I => \N__31091\
        );

    \I__6786\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31088\
        );

    \I__6785\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31082\
        );

    \I__6784\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31082\
        );

    \I__6783\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31079\
        );

    \I__6782\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31076\
        );

    \I__6781\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31073\
        );

    \I__6780\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31070\
        );

    \I__6779\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31067\
        );

    \I__6778\ : Span4Mux_v
    port map (
            O => \N__31104\,
            I => \N__31064\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__31101\,
            I => \N__31060\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__31098\,
            I => \N__31057\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__31095\,
            I => \N__31054\
        );

    \I__6774\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31051\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__31091\,
            I => \N__31048\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__31088\,
            I => \N__31045\
        );

    \I__6771\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31042\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__31082\,
            I => \N__31037\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__31079\,
            I => \N__31037\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__31076\,
            I => \N__31032\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__31032\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__31070\,
            I => \N__31027\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__31067\,
            I => \N__31027\
        );

    \I__6764\ : Span4Mux_h
    port map (
            O => \N__31064\,
            I => \N__31024\
        );

    \I__6763\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31021\
        );

    \I__6762\ : Span4Mux_v
    port map (
            O => \N__31060\,
            I => \N__31018\
        );

    \I__6761\ : Span4Mux_h
    port map (
            O => \N__31057\,
            I => \N__31011\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__31054\,
            I => \N__31011\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__31051\,
            I => \N__31011\
        );

    \I__6758\ : Span4Mux_v
    port map (
            O => \N__31048\,
            I => \N__31004\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__31045\,
            I => \N__31004\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__31042\,
            I => \N__31004\
        );

    \I__6755\ : Span4Mux_v
    port map (
            O => \N__31037\,
            I => \N__31001\
        );

    \I__6754\ : Span4Mux_h
    port map (
            O => \N__31032\,
            I => \N__30996\
        );

    \I__6753\ : Span4Mux_h
    port map (
            O => \N__31027\,
            I => \N__30996\
        );

    \I__6752\ : Span4Mux_h
    port map (
            O => \N__31024\,
            I => \N__30991\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__31021\,
            I => \N__30991\
        );

    \I__6750\ : Span4Mux_v
    port map (
            O => \N__31018\,
            I => \N__30988\
        );

    \I__6749\ : Span4Mux_v
    port map (
            O => \N__31011\,
            I => \N__30981\
        );

    \I__6748\ : Span4Mux_h
    port map (
            O => \N__31004\,
            I => \N__30981\
        );

    \I__6747\ : Span4Mux_v
    port map (
            O => \N__31001\,
            I => \N__30981\
        );

    \I__6746\ : Span4Mux_v
    port map (
            O => \N__30996\,
            I => \N__30978\
        );

    \I__6745\ : Odrv4
    port map (
            O => \N__30991\,
            I => \dataWriteZ0Z_6\
        );

    \I__6744\ : Odrv4
    port map (
            O => \N__30988\,
            I => \dataWriteZ0Z_6\
        );

    \I__6743\ : Odrv4
    port map (
            O => \N__30981\,
            I => \dataWriteZ0Z_6\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__30978\,
            I => \dataWriteZ0Z_6\
        );

    \I__6741\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__30966\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_6\
        );

    \I__6739\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30960\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__30960\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_8\
        );

    \I__6737\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30954\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__30954\,
            I => \PWMInstance2.PWMPulseWidthCountZ0Z_9\
        );

    \I__6735\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30948\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__30948\,
            I => \N__30944\
        );

    \I__6733\ : CascadeMux
    port map (
            O => \N__30947\,
            I => \N__30940\
        );

    \I__6732\ : Span4Mux_h
    port map (
            O => \N__30944\,
            I => \N__30937\
        );

    \I__6731\ : CascadeMux
    port map (
            O => \N__30943\,
            I => \N__30934\
        );

    \I__6730\ : InMux
    port map (
            O => \N__30940\,
            I => \N__30931\
        );

    \I__6729\ : Span4Mux_h
    port map (
            O => \N__30937\,
            I => \N__30928\
        );

    \I__6728\ : InMux
    port map (
            O => \N__30934\,
            I => \N__30925\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__30931\,
            I => \dataRead1_0\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__30928\,
            I => \dataRead1_0\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__30925\,
            I => \dataRead1_0\
        );

    \I__6724\ : CascadeMux
    port map (
            O => \N__30918\,
            I => \OutReg_0_5_i_m3_ns_1_0_cascade_\
        );

    \I__6723\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30912\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N__30909\
        );

    \I__6721\ : Span4Mux_h
    port map (
            O => \N__30909\,
            I => \N__30904\
        );

    \I__6720\ : CascadeMux
    port map (
            O => \N__30908\,
            I => \N__30901\
        );

    \I__6719\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30898\
        );

    \I__6718\ : Span4Mux_v
    port map (
            O => \N__30904\,
            I => \N__30895\
        );

    \I__6717\ : InMux
    port map (
            O => \N__30901\,
            I => \N__30892\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__30898\,
            I => \dataRead5_0\
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__30895\,
            I => \dataRead5_0\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__30892\,
            I => \dataRead5_0\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__30885\,
            I => \OutReg_ess_RNO_1Z0Z_0_cascade_\
        );

    \I__6712\ : InMux
    port map (
            O => \N__30882\,
            I => \N__30879\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__30879\,
            I => \N__30874\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__30878\,
            I => \N__30871\
        );

    \I__6709\ : InMux
    port map (
            O => \N__30877\,
            I => \N__30868\
        );

    \I__6708\ : Span4Mux_v
    port map (
            O => \N__30874\,
            I => \N__30865\
        );

    \I__6707\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30862\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__30868\,
            I => \N__30857\
        );

    \I__6705\ : Span4Mux_h
    port map (
            O => \N__30865\,
            I => \N__30857\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__30862\,
            I => \N__30854\
        );

    \I__6703\ : Odrv4
    port map (
            O => \N__30857\,
            I => \dataRead3_0\
        );

    \I__6702\ : Odrv12
    port map (
            O => \N__30854\,
            I => \dataRead3_0\
        );

    \I__6701\ : CascadeMux
    port map (
            O => \N__30849\,
            I => \N__30846\
        );

    \I__6700\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30842\
        );

    \I__6699\ : CascadeMux
    port map (
            O => \N__30845\,
            I => \N__30839\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__30842\,
            I => \N__30835\
        );

    \I__6697\ : InMux
    port map (
            O => \N__30839\,
            I => \N__30832\
        );

    \I__6696\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30829\
        );

    \I__6695\ : Span4Mux_v
    port map (
            O => \N__30835\,
            I => \N__30826\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__30832\,
            I => \N__30823\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__30829\,
            I => \N__30818\
        );

    \I__6692\ : Span4Mux_h
    port map (
            O => \N__30826\,
            I => \N__30818\
        );

    \I__6691\ : Span4Mux_h
    port map (
            O => \N__30823\,
            I => \N__30815\
        );

    \I__6690\ : Odrv4
    port map (
            O => \N__30818\,
            I => \dataRead2_0\
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__30815\,
            I => \dataRead2_0\
        );

    \I__6688\ : CascadeMux
    port map (
            O => \N__30810\,
            I => \N__30806\
        );

    \I__6687\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30803\
        );

    \I__6686\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30800\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__30803\,
            I => \N__30796\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__30800\,
            I => \N__30793\
        );

    \I__6683\ : InMux
    port map (
            O => \N__30799\,
            I => \N__30790\
        );

    \I__6682\ : Span4Mux_h
    port map (
            O => \N__30796\,
            I => \N__30785\
        );

    \I__6681\ : Span4Mux_h
    port map (
            O => \N__30793\,
            I => \N__30785\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__30790\,
            I => \dataRead6_0\
        );

    \I__6679\ : Odrv4
    port map (
            O => \N__30785\,
            I => \dataRead6_0\
        );

    \I__6678\ : CascadeMux
    port map (
            O => \N__30780\,
            I => \OutReg_0_4_i_m3_ns_1_0_cascade_\
        );

    \I__6677\ : InMux
    port map (
            O => \N__30777\,
            I => \N__30773\
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__30776\,
            I => \N__30770\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__30773\,
            I => \N__30766\
        );

    \I__6674\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30763\
        );

    \I__6673\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30760\
        );

    \I__6672\ : Span4Mux_h
    port map (
            O => \N__30766\,
            I => \N__30757\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__30763\,
            I => \N__30754\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__30760\,
            I => \dataRead7_0\
        );

    \I__6669\ : Odrv4
    port map (
            O => \N__30757\,
            I => \dataRead7_0\
        );

    \I__6668\ : Odrv12
    port map (
            O => \N__30754\,
            I => \dataRead7_0\
        );

    \I__6667\ : InMux
    port map (
            O => \N__30747\,
            I => \N__30744\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__30744\,
            I => \OutReg_ess_RNO_0Z0Z_0\
        );

    \I__6665\ : CascadeMux
    port map (
            O => \N__30741\,
            I => \N__30738\
        );

    \I__6664\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30735\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__30735\,
            I => \N__30732\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__30732\,
            I => \OutRegZ0Z_0\
        );

    \I__6661\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30726\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__30726\,
            I => \N__30723\
        );

    \I__6659\ : Span4Mux_h
    port map (
            O => \N__30723\,
            I => \N__30720\
        );

    \I__6658\ : Odrv4
    port map (
            O => \N__30720\,
            I => \OutReg_ess_RNO_0Z0Z_1\
        );

    \I__6657\ : InMux
    port map (
            O => \N__30717\,
            I => \N__30714\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__30714\,
            I => \OutRegZ0Z_1\
        );

    \I__6655\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30707\
        );

    \I__6654\ : InMux
    port map (
            O => \N__30710\,
            I => \N__30704\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__30707\,
            I => \N__30700\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__30704\,
            I => \N__30697\
        );

    \I__6651\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30694\
        );

    \I__6650\ : Span4Mux_v
    port map (
            O => \N__30700\,
            I => \N__30691\
        );

    \I__6649\ : Span4Mux_h
    port map (
            O => \N__30697\,
            I => \N__30688\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__30694\,
            I => \N__30685\
        );

    \I__6647\ : Span4Mux_h
    port map (
            O => \N__30691\,
            I => \N__30680\
        );

    \I__6646\ : Span4Mux_h
    port map (
            O => \N__30688\,
            I => \N__30680\
        );

    \I__6645\ : Odrv12
    port map (
            O => \N__30685\,
            I => \dataRead2_8\
        );

    \I__6644\ : Odrv4
    port map (
            O => \N__30680\,
            I => \dataRead2_8\
        );

    \I__6643\ : CascadeMux
    port map (
            O => \N__30675\,
            I => \N__30672\
        );

    \I__6642\ : InMux
    port map (
            O => \N__30672\,
            I => \N__30669\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__30669\,
            I => \N__30665\
        );

    \I__6640\ : InMux
    port map (
            O => \N__30668\,
            I => \N__30662\
        );

    \I__6639\ : Span4Mux_h
    port map (
            O => \N__30665\,
            I => \N__30658\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__30662\,
            I => \N__30655\
        );

    \I__6637\ : InMux
    port map (
            O => \N__30661\,
            I => \N__30652\
        );

    \I__6636\ : Span4Mux_h
    port map (
            O => \N__30658\,
            I => \N__30649\
        );

    \I__6635\ : Odrv4
    port map (
            O => \N__30655\,
            I => \dataRead3_8\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__30652\,
            I => \dataRead3_8\
        );

    \I__6633\ : Odrv4
    port map (
            O => \N__30649\,
            I => \dataRead3_8\
        );

    \I__6632\ : CascadeMux
    port map (
            O => \N__30642\,
            I => \N__30639\
        );

    \I__6631\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30635\
        );

    \I__6630\ : InMux
    port map (
            O => \N__30638\,
            I => \N__30631\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__30635\,
            I => \N__30628\
        );

    \I__6628\ : InMux
    port map (
            O => \N__30634\,
            I => \N__30625\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__30631\,
            I => \N__30622\
        );

    \I__6626\ : Span4Mux_h
    port map (
            O => \N__30628\,
            I => \N__30616\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__30625\,
            I => \N__30616\
        );

    \I__6624\ : Span4Mux_h
    port map (
            O => \N__30622\,
            I => \N__30613\
        );

    \I__6623\ : InMux
    port map (
            O => \N__30621\,
            I => \N__30610\
        );

    \I__6622\ : Span4Mux_h
    port map (
            O => \N__30616\,
            I => \N__30607\
        );

    \I__6621\ : Odrv4
    port map (
            O => \N__30613\,
            I => \data_receivedZ0Z_3\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__30610\,
            I => \data_receivedZ0Z_3\
        );

    \I__6619\ : Odrv4
    port map (
            O => \N__30607\,
            I => \data_receivedZ0Z_3\
        );

    \I__6618\ : CascadeMux
    port map (
            O => \N__30600\,
            I => \data_received_esr_RNI7L871Z0Z_3_cascade_\
        );

    \I__6617\ : InMux
    port map (
            O => \N__30597\,
            I => \QuadInstance0.un1_Quad_cry_13\
        );

    \I__6616\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30591\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__30591\,
            I => \N__30588\
        );

    \I__6614\ : Odrv4
    port map (
            O => \N__30588\,
            I => \QuadInstance0.un1_Quad_axb_15\
        );

    \I__6613\ : InMux
    port map (
            O => \N__30585\,
            I => \QuadInstance0.un1_Quad_cry_14\
        );

    \I__6612\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30576\
        );

    \I__6611\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30576\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__30576\,
            I => \N__30573\
        );

    \I__6609\ : Odrv4
    port map (
            O => \N__30573\,
            I => \dataRead0_15\
        );

    \I__6608\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30565\
        );

    \I__6607\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30562\
        );

    \I__6606\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30559\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__30565\,
            I => \N__30556\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__30562\,
            I => \N__30551\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30551\
        );

    \I__6602\ : Span4Mux_v
    port map (
            O => \N__30556\,
            I => \N__30548\
        );

    \I__6601\ : Span4Mux_h
    port map (
            O => \N__30551\,
            I => \N__30545\
        );

    \I__6600\ : Sp12to4
    port map (
            O => \N__30548\,
            I => \N__30542\
        );

    \I__6599\ : Span4Mux_h
    port map (
            O => \N__30545\,
            I => \N__30539\
        );

    \I__6598\ : Odrv12
    port map (
            O => \N__30542\,
            I => \dataRead1_2\
        );

    \I__6597\ : Odrv4
    port map (
            O => \N__30539\,
            I => \dataRead1_2\
        );

    \I__6596\ : CascadeMux
    port map (
            O => \N__30534\,
            I => \N__30531\
        );

    \I__6595\ : InMux
    port map (
            O => \N__30531\,
            I => \N__30527\
        );

    \I__6594\ : InMux
    port map (
            O => \N__30530\,
            I => \N__30523\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__30527\,
            I => \N__30520\
        );

    \I__6592\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30517\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__30523\,
            I => \N__30514\
        );

    \I__6590\ : Span4Mux_h
    port map (
            O => \N__30520\,
            I => \N__30511\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__30517\,
            I => \N__30508\
        );

    \I__6588\ : Span4Mux_h
    port map (
            O => \N__30514\,
            I => \N__30505\
        );

    \I__6587\ : Span4Mux_h
    port map (
            O => \N__30511\,
            I => \N__30502\
        );

    \I__6586\ : Span4Mux_v
    port map (
            O => \N__30508\,
            I => \N__30499\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__30505\,
            I => \dataRead5_2\
        );

    \I__6584\ : Odrv4
    port map (
            O => \N__30502\,
            I => \dataRead5_2\
        );

    \I__6583\ : Odrv4
    port map (
            O => \N__30499\,
            I => \dataRead5_2\
        );

    \I__6582\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__30489\,
            I => \N__30486\
        );

    \I__6580\ : Span4Mux_v
    port map (
            O => \N__30486\,
            I => \N__30483\
        );

    \I__6579\ : Odrv4
    port map (
            O => \N__30483\,
            I => \OutReg_0_5_i_m3_ns_1_2\
        );

    \I__6578\ : CascadeMux
    port map (
            O => \N__30480\,
            I => \OutReg_esr_RNO_2Z0Z_2_cascade_\
        );

    \I__6577\ : CascadeMux
    port map (
            O => \N__30477\,
            I => \OutReg_esr_RNO_0Z0Z_2_cascade_\
        );

    \I__6576\ : InMux
    port map (
            O => \N__30474\,
            I => \N__30471\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__30471\,
            I => \N__30468\
        );

    \I__6574\ : Odrv4
    port map (
            O => \N__30468\,
            I => \OutRegZ0Z_2\
        );

    \I__6573\ : InMux
    port map (
            O => \N__30465\,
            I => \N__30462\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__30462\,
            I => \N__30457\
        );

    \I__6571\ : InMux
    port map (
            O => \N__30461\,
            I => \N__30454\
        );

    \I__6570\ : InMux
    port map (
            O => \N__30460\,
            I => \N__30451\
        );

    \I__6569\ : Span4Mux_v
    port map (
            O => \N__30457\,
            I => \N__30446\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__30454\,
            I => \N__30446\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__30451\,
            I => \N__30443\
        );

    \I__6566\ : Span4Mux_h
    port map (
            O => \N__30446\,
            I => \N__30440\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__30443\,
            I => \N__30437\
        );

    \I__6564\ : Span4Mux_h
    port map (
            O => \N__30440\,
            I => \N__30434\
        );

    \I__6563\ : Span4Mux_h
    port map (
            O => \N__30437\,
            I => \N__30431\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__30434\,
            I => \dataRead2_2\
        );

    \I__6561\ : Odrv4
    port map (
            O => \N__30431\,
            I => \dataRead2_2\
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__30426\,
            I => \N__30423\
        );

    \I__6559\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30419\
        );

    \I__6558\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30415\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__30419\,
            I => \N__30412\
        );

    \I__6556\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30409\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__30415\,
            I => \N__30406\
        );

    \I__6554\ : Span4Mux_h
    port map (
            O => \N__30412\,
            I => \N__30403\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__30409\,
            I => \N__30400\
        );

    \I__6552\ : Sp12to4
    port map (
            O => \N__30406\,
            I => \N__30397\
        );

    \I__6551\ : Span4Mux_v
    port map (
            O => \N__30403\,
            I => \N__30392\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__30400\,
            I => \N__30392\
        );

    \I__6549\ : Odrv12
    port map (
            O => \N__30397\,
            I => \dataRead3_2\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__30392\,
            I => \dataRead3_2\
        );

    \I__6547\ : InMux
    port map (
            O => \N__30387\,
            I => \N__30383\
        );

    \I__6546\ : InMux
    port map (
            O => \N__30386\,
            I => \N__30380\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__30383\,
            I => \N__30376\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__30380\,
            I => \N__30373\
        );

    \I__6543\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30370\
        );

    \I__6542\ : Span4Mux_v
    port map (
            O => \N__30376\,
            I => \N__30367\
        );

    \I__6541\ : Span4Mux_v
    port map (
            O => \N__30373\,
            I => \N__30362\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__30370\,
            I => \N__30362\
        );

    \I__6539\ : Span4Mux_h
    port map (
            O => \N__30367\,
            I => \N__30357\
        );

    \I__6538\ : Span4Mux_v
    port map (
            O => \N__30362\,
            I => \N__30357\
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__30357\,
            I => \dataRead7_2\
        );

    \I__6536\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30350\
        );

    \I__6535\ : InMux
    port map (
            O => \N__30353\,
            I => \N__30347\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__30350\,
            I => \N__30341\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30341\
        );

    \I__6532\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30338\
        );

    \I__6531\ : Span12Mux_h
    port map (
            O => \N__30341\,
            I => \N__30335\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__30338\,
            I => \N__30332\
        );

    \I__6529\ : Odrv12
    port map (
            O => \N__30335\,
            I => \dataRead6_2\
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__30332\,
            I => \dataRead6_2\
        );

    \I__6527\ : CascadeMux
    port map (
            O => \N__30327\,
            I => \OutReg_0_4_i_m3_ns_1_2_cascade_\
        );

    \I__6526\ : InMux
    port map (
            O => \N__30324\,
            I => \N__30321\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__30321\,
            I => \OutReg_esr_RNO_1Z0Z_2\
        );

    \I__6524\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30314\
        );

    \I__6523\ : CascadeMux
    port map (
            O => \N__30317\,
            I => \N__30311\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__30314\,
            I => \N__30308\
        );

    \I__6521\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30305\
        );

    \I__6520\ : Span4Mux_v
    port map (
            O => \N__30308\,
            I => \N__30300\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__30305\,
            I => \N__30300\
        );

    \I__6518\ : Span4Mux_h
    port map (
            O => \N__30300\,
            I => \N__30296\
        );

    \I__6517\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30293\
        );

    \I__6516\ : Span4Mux_h
    port map (
            O => \N__30296\,
            I => \N__30290\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__30293\,
            I => \dataRead0_0\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__30290\,
            I => \dataRead0_0\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__30285\,
            I => \N__30281\
        );

    \I__6512\ : CascadeMux
    port map (
            O => \N__30284\,
            I => \N__30278\
        );

    \I__6511\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30275\
        );

    \I__6510\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30272\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__30275\,
            I => \N__30269\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__30272\,
            I => \N__30265\
        );

    \I__6507\ : Span4Mux_v
    port map (
            O => \N__30269\,
            I => \N__30262\
        );

    \I__6506\ : InMux
    port map (
            O => \N__30268\,
            I => \N__30259\
        );

    \I__6505\ : Span4Mux_s2_v
    port map (
            O => \N__30265\,
            I => \N__30256\
        );

    \I__6504\ : Span4Mux_h
    port map (
            O => \N__30262\,
            I => \N__30253\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__30259\,
            I => \N__30248\
        );

    \I__6502\ : Span4Mux_h
    port map (
            O => \N__30256\,
            I => \N__30248\
        );

    \I__6501\ : Odrv4
    port map (
            O => \N__30253\,
            I => \dataRead4_0\
        );

    \I__6500\ : Odrv4
    port map (
            O => \N__30248\,
            I => \dataRead4_0\
        );

    \I__6499\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__30240\,
            I => \N__30237\
        );

    \I__6497\ : Span4Mux_h
    port map (
            O => \N__30237\,
            I => \N__30234\
        );

    \I__6496\ : Odrv4
    port map (
            O => \N__30234\,
            I => \QuadInstance0.Quad_RNO_0_0_6\
        );

    \I__6495\ : InMux
    port map (
            O => \N__30231\,
            I => \QuadInstance0.un1_Quad_cry_5\
        );

    \I__6494\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30223\
        );

    \I__6493\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30218\
        );

    \I__6492\ : InMux
    port map (
            O => \N__30226\,
            I => \N__30218\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__30223\,
            I => \dataRead0_7\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__30218\,
            I => \dataRead0_7\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__30213\,
            I => \N__30210\
        );

    \I__6488\ : InMux
    port map (
            O => \N__30210\,
            I => \N__30207\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__30207\,
            I => \QuadInstance0.Quad_RNIMKBH1Z0Z_7\
        );

    \I__6486\ : InMux
    port map (
            O => \N__30204\,
            I => \N__30201\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__30201\,
            I => \QuadInstance0.Quad_RNO_0_0_7\
        );

    \I__6484\ : InMux
    port map (
            O => \N__30198\,
            I => \QuadInstance0.un1_Quad_cry_6\
        );

    \I__6483\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30190\
        );

    \I__6482\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30185\
        );

    \I__6481\ : InMux
    port map (
            O => \N__30193\,
            I => \N__30185\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__30190\,
            I => \dataRead0_8\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__30185\,
            I => \dataRead0_8\
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__30180\,
            I => \N__30177\
        );

    \I__6477\ : InMux
    port map (
            O => \N__30177\,
            I => \N__30174\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__30174\,
            I => \QuadInstance0.Quad_RNINLBH1Z0Z_8\
        );

    \I__6475\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30168\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__30168\,
            I => \QuadInstance0.Quad_RNO_0_0_8\
        );

    \I__6473\ : InMux
    port map (
            O => \N__30165\,
            I => \bfn_17_7_0_\
        );

    \I__6472\ : InMux
    port map (
            O => \N__30162\,
            I => \N__30158\
        );

    \I__6471\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30154\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__30158\,
            I => \N__30151\
        );

    \I__6469\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30148\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__30154\,
            I => \N__30145\
        );

    \I__6467\ : Span4Mux_v
    port map (
            O => \N__30151\,
            I => \N__30140\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__30148\,
            I => \N__30140\
        );

    \I__6465\ : Span4Mux_v
    port map (
            O => \N__30145\,
            I => \N__30137\
        );

    \I__6464\ : Span4Mux_h
    port map (
            O => \N__30140\,
            I => \N__30134\
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__30137\,
            I => \dataRead0_9\
        );

    \I__6462\ : Odrv4
    port map (
            O => \N__30134\,
            I => \dataRead0_9\
        );

    \I__6461\ : CascadeMux
    port map (
            O => \N__30129\,
            I => \N__30126\
        );

    \I__6460\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30123\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__30123\,
            I => \N__30120\
        );

    \I__6458\ : Odrv4
    port map (
            O => \N__30120\,
            I => \QuadInstance0.Quad_RNIOMBH1Z0Z_9\
        );

    \I__6457\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__30114\,
            I => \N__30111\
        );

    \I__6455\ : Span4Mux_h
    port map (
            O => \N__30111\,
            I => \N__30108\
        );

    \I__6454\ : Odrv4
    port map (
            O => \N__30108\,
            I => \QuadInstance0.Quad_RNO_0_0_9\
        );

    \I__6453\ : InMux
    port map (
            O => \N__30105\,
            I => \QuadInstance0.un1_Quad_cry_8\
        );

    \I__6452\ : InMux
    port map (
            O => \N__30102\,
            I => \QuadInstance0.un1_Quad_cry_9\
        );

    \I__6451\ : InMux
    port map (
            O => \N__30099\,
            I => \N__30094\
        );

    \I__6450\ : InMux
    port map (
            O => \N__30098\,
            I => \N__30091\
        );

    \I__6449\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30088\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__30094\,
            I => \N__30083\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__30091\,
            I => \N__30083\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__30088\,
            I => \N__30080\
        );

    \I__6445\ : Odrv12
    port map (
            O => \N__30083\,
            I => \dataRead0_11\
        );

    \I__6444\ : Odrv12
    port map (
            O => \N__30080\,
            I => \dataRead0_11\
        );

    \I__6443\ : CascadeMux
    port map (
            O => \N__30075\,
            I => \N__30072\
        );

    \I__6442\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30069\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__30069\,
            I => \QuadInstance0.Quad_RNI1M8Q1Z0Z_11\
        );

    \I__6440\ : InMux
    port map (
            O => \N__30066\,
            I => \N__30063\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__30063\,
            I => \N__30060\
        );

    \I__6438\ : Odrv12
    port map (
            O => \N__30060\,
            I => \QuadInstance0.Quad_RNO_0_0_11\
        );

    \I__6437\ : InMux
    port map (
            O => \N__30057\,
            I => \QuadInstance0.un1_Quad_cry_10\
        );

    \I__6436\ : InMux
    port map (
            O => \N__30054\,
            I => \N__30050\
        );

    \I__6435\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30046\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__30050\,
            I => \N__30043\
        );

    \I__6433\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30040\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__30046\,
            I => \dataRead0_12\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__30043\,
            I => \dataRead0_12\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__30040\,
            I => \dataRead0_12\
        );

    \I__6429\ : CascadeMux
    port map (
            O => \N__30033\,
            I => \N__30030\
        );

    \I__6428\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30027\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__30027\,
            I => \QuadInstance0.Quad_RNI2N8Q1Z0Z_12\
        );

    \I__6426\ : InMux
    port map (
            O => \N__30024\,
            I => \N__30021\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__30021\,
            I => \QuadInstance0.Quad_RNO_0_0_12\
        );

    \I__6424\ : InMux
    port map (
            O => \N__30018\,
            I => \QuadInstance0.un1_Quad_cry_11\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__30015\,
            I => \N__30010\
        );

    \I__6422\ : InMux
    port map (
            O => \N__30014\,
            I => \N__30007\
        );

    \I__6421\ : InMux
    port map (
            O => \N__30013\,
            I => \N__30002\
        );

    \I__6420\ : InMux
    port map (
            O => \N__30010\,
            I => \N__30002\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__30007\,
            I => \dataRead0_13\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__30002\,
            I => \dataRead0_13\
        );

    \I__6417\ : CascadeMux
    port map (
            O => \N__29997\,
            I => \N__29994\
        );

    \I__6416\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29991\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__29991\,
            I => \QuadInstance0.Quad_RNI3O8Q1Z0Z_13\
        );

    \I__6414\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29985\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__29985\,
            I => \QuadInstance0.Quad_RNO_0_0_13\
        );

    \I__6412\ : InMux
    port map (
            O => \N__29982\,
            I => \QuadInstance0.un1_Quad_cry_12\
        );

    \I__6411\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29976\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__29976\,
            I => \N__29973\
        );

    \I__6409\ : Odrv4
    port map (
            O => \N__29973\,
            I => \QuadInstance4.Quad_RNO_0_4_14\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__29970\,
            I => \N__29966\
        );

    \I__6407\ : CascadeMux
    port map (
            O => \N__29969\,
            I => \N__29962\
        );

    \I__6406\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29959\
        );

    \I__6405\ : CascadeMux
    port map (
            O => \N__29965\,
            I => \N__29956\
        );

    \I__6404\ : InMux
    port map (
            O => \N__29962\,
            I => \N__29953\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__29959\,
            I => \N__29950\
        );

    \I__6402\ : InMux
    port map (
            O => \N__29956\,
            I => \N__29947\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__29953\,
            I => \N__29944\
        );

    \I__6400\ : Span4Mux_v
    port map (
            O => \N__29950\,
            I => \N__29941\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__29947\,
            I => \dataRead4_14\
        );

    \I__6398\ : Odrv12
    port map (
            O => \N__29944\,
            I => \dataRead4_14\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__29941\,
            I => \dataRead4_14\
        );

    \I__6396\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29931\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__29931\,
            I => \N__29928\
        );

    \I__6394\ : Span4Mux_v
    port map (
            O => \N__29928\,
            I => \N__29925\
        );

    \I__6393\ : Sp12to4
    port map (
            O => \N__29925\,
            I => \N__29922\
        );

    \I__6392\ : Odrv12
    port map (
            O => \N__29922\,
            I => \QuadInstance0.delayedCh_BZ0Z_0\
        );

    \I__6391\ : InMux
    port map (
            O => \N__29919\,
            I => \N__29916\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__29916\,
            I => \N__29913\
        );

    \I__6389\ : Span4Mux_h
    port map (
            O => \N__29913\,
            I => \N__29910\
        );

    \I__6388\ : Odrv4
    port map (
            O => \N__29910\,
            I => \QuadInstance4.delayedCh_BZ0Z_0\
        );

    \I__6387\ : CascadeMux
    port map (
            O => \N__29907\,
            I => \N__29903\
        );

    \I__6386\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29900\
        );

    \I__6385\ : InMux
    port map (
            O => \N__29903\,
            I => \N__29897\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__29900\,
            I => \QuadInstance4.delayedCh_BZ0Z_1\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__29897\,
            I => \QuadInstance4.delayedCh_BZ0Z_1\
        );

    \I__6382\ : InMux
    port map (
            O => \N__29892\,
            I => \N__29889\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__29889\,
            I => \N__29886\
        );

    \I__6380\ : Span4Mux_h
    port map (
            O => \N__29886\,
            I => \N__29883\
        );

    \I__6379\ : Odrv4
    port map (
            O => \N__29883\,
            I => \QuadInstance0.Quad_RNO_0Z0Z_1\
        );

    \I__6378\ : InMux
    port map (
            O => \N__29880\,
            I => \QuadInstance0.un1_Quad_cry_0\
        );

    \I__6377\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29874\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__29874\,
            I => \N__29871\
        );

    \I__6375\ : Odrv4
    port map (
            O => \N__29871\,
            I => \QuadInstance0.Quad_RNO_0_0_2\
        );

    \I__6374\ : InMux
    port map (
            O => \N__29868\,
            I => \QuadInstance0.un1_Quad_cry_1\
        );

    \I__6373\ : InMux
    port map (
            O => \N__29865\,
            I => \N__29862\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__29862\,
            I => \N__29859\
        );

    \I__6371\ : Span4Mux_h
    port map (
            O => \N__29859\,
            I => \N__29856\
        );

    \I__6370\ : Span4Mux_h
    port map (
            O => \N__29856\,
            I => \N__29853\
        );

    \I__6369\ : Odrv4
    port map (
            O => \N__29853\,
            I => \QuadInstance0.Quad_RNO_0_0_3\
        );

    \I__6368\ : InMux
    port map (
            O => \N__29850\,
            I => \QuadInstance0.un1_Quad_cry_2\
        );

    \I__6367\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29844\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__29844\,
            I => \N__29841\
        );

    \I__6365\ : Span4Mux_h
    port map (
            O => \N__29841\,
            I => \N__29838\
        );

    \I__6364\ : Odrv4
    port map (
            O => \N__29838\,
            I => \QuadInstance0.Quad_RNO_0_0_4\
        );

    \I__6363\ : InMux
    port map (
            O => \N__29835\,
            I => \QuadInstance0.un1_Quad_cry_3\
        );

    \I__6362\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29829\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__29829\,
            I => \N__29826\
        );

    \I__6360\ : Odrv4
    port map (
            O => \N__29826\,
            I => \QuadInstance0.Quad_RNO_0_0_5\
        );

    \I__6359\ : InMux
    port map (
            O => \N__29823\,
            I => \QuadInstance0.un1_Quad_cry_4\
        );

    \I__6358\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29817\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__29817\,
            I => \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_2\
        );

    \I__6356\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29811\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__29811\,
            I => \N__29808\
        );

    \I__6354\ : Odrv4
    port map (
            O => \N__29808\,
            I => \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_2\
        );

    \I__6353\ : InMux
    port map (
            O => \N__29805\,
            I => \N__29802\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__29802\,
            I => \N__29799\
        );

    \I__6351\ : Odrv4
    port map (
            O => \N__29799\,
            I => \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_2\
        );

    \I__6350\ : InMux
    port map (
            O => \N__29796\,
            I => \N__29793\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__6348\ : Odrv4
    port map (
            O => \N__29790\,
            I => \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_2\
        );

    \I__6347\ : InMux
    port map (
            O => \N__29787\,
            I => \N__29784\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__29784\,
            I => \N__29781\
        );

    \I__6345\ : Span4Mux_v
    port map (
            O => \N__29781\,
            I => \N__29778\
        );

    \I__6344\ : Odrv4
    port map (
            O => \N__29778\,
            I => \PWMInstance3.un1_periodCounter12_1_0_a2_0\
        );

    \I__6343\ : CascadeMux
    port map (
            O => \N__29775\,
            I => \N__29772\
        );

    \I__6342\ : InMux
    port map (
            O => \N__29772\,
            I => \N__29768\
        );

    \I__6341\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29761\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__29768\,
            I => \N__29758\
        );

    \I__6339\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29753\
        );

    \I__6338\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29753\
        );

    \I__6337\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29750\
        );

    \I__6336\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29747\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__29761\,
            I => \N__29744\
        );

    \I__6334\ : Span4Mux_h
    port map (
            O => \N__29758\,
            I => \N__29741\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__29753\,
            I => \PWMInstance3.out_0_sqmuxa\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__29750\,
            I => \PWMInstance3.out_0_sqmuxa\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__29747\,
            I => \PWMInstance3.out_0_sqmuxa\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__29744\,
            I => \PWMInstance3.out_0_sqmuxa\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__29741\,
            I => \PWMInstance3.out_0_sqmuxa\
        );

    \I__6328\ : InMux
    port map (
            O => \N__29730\,
            I => \bfn_16_16_0_\
        );

    \I__6327\ : IoInMux
    port map (
            O => \N__29727\,
            I => \N__29724\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__29724\,
            I => \N__29721\
        );

    \I__6325\ : Span4Mux_s0_v
    port map (
            O => \N__29721\,
            I => \N__29718\
        );

    \I__6324\ : Span4Mux_v
    port map (
            O => \N__29718\,
            I => \N__29714\
        );

    \I__6323\ : InMux
    port map (
            O => \N__29717\,
            I => \N__29711\
        );

    \I__6322\ : Odrv4
    port map (
            O => \N__29714\,
            I => \PWM3_c\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__29711\,
            I => \PWM3_c\
        );

    \I__6320\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29703\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__29703\,
            I => \N__29700\
        );

    \I__6318\ : IoSpan4Mux
    port map (
            O => \N__29700\,
            I => \N__29697\
        );

    \I__6317\ : Odrv4
    port map (
            O => \N__29697\,
            I => \ch7_A_c\
        );

    \I__6316\ : InMux
    port map (
            O => \N__29694\,
            I => \N__29691\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__29691\,
            I => \N__29688\
        );

    \I__6314\ : Span4Mux_h
    port map (
            O => \N__29688\,
            I => \N__29685\
        );

    \I__6313\ : Span4Mux_v
    port map (
            O => \N__29685\,
            I => \N__29682\
        );

    \I__6312\ : Span4Mux_h
    port map (
            O => \N__29682\,
            I => \N__29679\
        );

    \I__6311\ : Odrv4
    port map (
            O => \N__29679\,
            I => \QuadInstance7.delayedCh_AZ0Z_0\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__29676\,
            I => \N__29673\
        );

    \I__6309\ : InMux
    port map (
            O => \N__29673\,
            I => \N__29670\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__29670\,
            I => \N__29667\
        );

    \I__6307\ : Odrv4
    port map (
            O => \N__29667\,
            I => \QuadInstance4.Quad_RNO_0_4_10\
        );

    \I__6306\ : InMux
    port map (
            O => \N__29664\,
            I => \N__29653\
        );

    \I__6305\ : InMux
    port map (
            O => \N__29663\,
            I => \N__29653\
        );

    \I__6304\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29649\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29644\
        );

    \I__6302\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29644\
        );

    \I__6301\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29637\
        );

    \I__6300\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29637\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__29653\,
            I => \N__29634\
        );

    \I__6298\ : CascadeMux
    port map (
            O => \N__29652\,
            I => \N__29630\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__29649\,
            I => \N__29625\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__29644\,
            I => \N__29615\
        );

    \I__6295\ : InMux
    port map (
            O => \N__29643\,
            I => \N__29610\
        );

    \I__6294\ : InMux
    port map (
            O => \N__29642\,
            I => \N__29610\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__29637\,
            I => \N__29605\
        );

    \I__6292\ : Span4Mux_h
    port map (
            O => \N__29634\,
            I => \N__29605\
        );

    \I__6291\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29591\
        );

    \I__6290\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29591\
        );

    \I__6289\ : InMux
    port map (
            O => \N__29629\,
            I => \N__29591\
        );

    \I__6288\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29584\
        );

    \I__6287\ : Span4Mux_h
    port map (
            O => \N__29625\,
            I => \N__29581\
        );

    \I__6286\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29572\
        );

    \I__6285\ : InMux
    port map (
            O => \N__29623\,
            I => \N__29572\
        );

    \I__6284\ : InMux
    port map (
            O => \N__29622\,
            I => \N__29572\
        );

    \I__6283\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29572\
        );

    \I__6282\ : InMux
    port map (
            O => \N__29620\,
            I => \N__29569\
        );

    \I__6281\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29564\
        );

    \I__6280\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29564\
        );

    \I__6279\ : Span4Mux_v
    port map (
            O => \N__29615\,
            I => \N__29561\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__29610\,
            I => \N__29556\
        );

    \I__6277\ : Span4Mux_h
    port map (
            O => \N__29605\,
            I => \N__29556\
        );

    \I__6276\ : InMux
    port map (
            O => \N__29604\,
            I => \N__29545\
        );

    \I__6275\ : InMux
    port map (
            O => \N__29603\,
            I => \N__29545\
        );

    \I__6274\ : InMux
    port map (
            O => \N__29602\,
            I => \N__29545\
        );

    \I__6273\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29545\
        );

    \I__6272\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29545\
        );

    \I__6271\ : InMux
    port map (
            O => \N__29599\,
            I => \N__29540\
        );

    \I__6270\ : InMux
    port map (
            O => \N__29598\,
            I => \N__29540\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__29591\,
            I => \N__29537\
        );

    \I__6268\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29528\
        );

    \I__6267\ : InMux
    port map (
            O => \N__29589\,
            I => \N__29528\
        );

    \I__6266\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29528\
        );

    \I__6265\ : InMux
    port map (
            O => \N__29587\,
            I => \N__29528\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__29584\,
            I => \N__29521\
        );

    \I__6263\ : Span4Mux_h
    port map (
            O => \N__29581\,
            I => \N__29521\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__29572\,
            I => \N__29521\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__29569\,
            I => \quadWriteZ0Z_4\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__29564\,
            I => \quadWriteZ0Z_4\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__29561\,
            I => \quadWriteZ0Z_4\
        );

    \I__6258\ : Odrv4
    port map (
            O => \N__29556\,
            I => \quadWriteZ0Z_4\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__29545\,
            I => \quadWriteZ0Z_4\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__29540\,
            I => \quadWriteZ0Z_4\
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__29537\,
            I => \quadWriteZ0Z_4\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__29528\,
            I => \quadWriteZ0Z_4\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__29521\,
            I => \quadWriteZ0Z_4\
        );

    \I__6252\ : CascadeMux
    port map (
            O => \N__29502\,
            I => \N__29498\
        );

    \I__6251\ : InMux
    port map (
            O => \N__29501\,
            I => \N__29494\
        );

    \I__6250\ : InMux
    port map (
            O => \N__29498\,
            I => \N__29491\
        );

    \I__6249\ : InMux
    port map (
            O => \N__29497\,
            I => \N__29488\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__29494\,
            I => \PWMInstance3.periodCounterZ0Z_7\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__29491\,
            I => \PWMInstance3.periodCounterZ0Z_7\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__29488\,
            I => \PWMInstance3.periodCounterZ0Z_7\
        );

    \I__6245\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29476\
        );

    \I__6244\ : InMux
    port map (
            O => \N__29480\,
            I => \N__29471\
        );

    \I__6243\ : InMux
    port map (
            O => \N__29479\,
            I => \N__29471\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__29476\,
            I => \PWMInstance3.periodCounterZ0Z_6\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__29471\,
            I => \PWMInstance3.periodCounterZ0Z_6\
        );

    \I__6240\ : InMux
    port map (
            O => \N__29466\,
            I => \N__29463\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__29463\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_6\
        );

    \I__6238\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__29457\,
            I => \N__29453\
        );

    \I__6236\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29445\
        );

    \I__6235\ : Span4Mux_v
    port map (
            O => \N__29453\,
            I => \N__29440\
        );

    \I__6234\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29431\
        );

    \I__6233\ : InMux
    port map (
            O => \N__29451\,
            I => \N__29431\
        );

    \I__6232\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29431\
        );

    \I__6231\ : InMux
    port map (
            O => \N__29449\,
            I => \N__29431\
        );

    \I__6230\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29428\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__29445\,
            I => \N__29422\
        );

    \I__6228\ : InMux
    port map (
            O => \N__29444\,
            I => \N__29419\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__29443\,
            I => \N__29414\
        );

    \I__6226\ : Span4Mux_h
    port map (
            O => \N__29440\,
            I => \N__29406\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__29431\,
            I => \N__29406\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__29428\,
            I => \N__29406\
        );

    \I__6223\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29401\
        );

    \I__6222\ : InMux
    port map (
            O => \N__29426\,
            I => \N__29401\
        );

    \I__6221\ : InMux
    port map (
            O => \N__29425\,
            I => \N__29398\
        );

    \I__6220\ : Span4Mux_h
    port map (
            O => \N__29422\,
            I => \N__29393\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__29419\,
            I => \N__29393\
        );

    \I__6218\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29389\
        );

    \I__6217\ : InMux
    port map (
            O => \N__29417\,
            I => \N__29386\
        );

    \I__6216\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29383\
        );

    \I__6215\ : InMux
    port map (
            O => \N__29413\,
            I => \N__29380\
        );

    \I__6214\ : Span4Mux_h
    port map (
            O => \N__29406\,
            I => \N__29375\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__29401\,
            I => \N__29375\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__29398\,
            I => \N__29372\
        );

    \I__6211\ : Span4Mux_h
    port map (
            O => \N__29393\,
            I => \N__29369\
        );

    \I__6210\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29366\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__29389\,
            I => \N__29363\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__29386\,
            I => \N__29358\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__29383\,
            I => \N__29358\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__29380\,
            I => \N__29355\
        );

    \I__6205\ : Span4Mux_h
    port map (
            O => \N__29375\,
            I => \N__29352\
        );

    \I__6204\ : Span4Mux_h
    port map (
            O => \N__29372\,
            I => \N__29349\
        );

    \I__6203\ : Span4Mux_v
    port map (
            O => \N__29369\,
            I => \N__29344\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__29366\,
            I => \N__29344\
        );

    \I__6201\ : Span12Mux_s11_h
    port map (
            O => \N__29363\,
            I => \N__29339\
        );

    \I__6200\ : Span12Mux_h
    port map (
            O => \N__29358\,
            I => \N__29339\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__29355\,
            I => \N__29334\
        );

    \I__6198\ : Span4Mux_v
    port map (
            O => \N__29352\,
            I => \N__29334\
        );

    \I__6197\ : Odrv4
    port map (
            O => \N__29349\,
            I => \dataWriteZ0Z_7\
        );

    \I__6196\ : Odrv4
    port map (
            O => \N__29344\,
            I => \dataWriteZ0Z_7\
        );

    \I__6195\ : Odrv12
    port map (
            O => \N__29339\,
            I => \dataWriteZ0Z_7\
        );

    \I__6194\ : Odrv4
    port map (
            O => \N__29334\,
            I => \dataWriteZ0Z_7\
        );

    \I__6193\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29322\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__29322\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_7\
        );

    \I__6191\ : CEMux
    port map (
            O => \N__29319\,
            I => \N__29315\
        );

    \I__6190\ : CEMux
    port map (
            O => \N__29318\,
            I => \N__29312\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__29315\,
            I => \N__29309\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__29312\,
            I => \N__29305\
        );

    \I__6187\ : Span4Mux_v
    port map (
            O => \N__29309\,
            I => \N__29302\
        );

    \I__6186\ : CEMux
    port map (
            O => \N__29308\,
            I => \N__29299\
        );

    \I__6185\ : Span4Mux_v
    port map (
            O => \N__29305\,
            I => \N__29291\
        );

    \I__6184\ : Span4Mux_v
    port map (
            O => \N__29302\,
            I => \N__29291\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__29299\,
            I => \N__29291\
        );

    \I__6182\ : CEMux
    port map (
            O => \N__29298\,
            I => \N__29287\
        );

    \I__6181\ : Span4Mux_v
    port map (
            O => \N__29291\,
            I => \N__29284\
        );

    \I__6180\ : CEMux
    port map (
            O => \N__29290\,
            I => \N__29281\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__29287\,
            I => \PWMInstance3.pwmWrite_0_3\
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__29284\,
            I => \PWMInstance3.pwmWrite_0_3\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__29281\,
            I => \PWMInstance3.pwmWrite_0_3\
        );

    \I__6176\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29271\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__29271\,
            I => \N__29268\
        );

    \I__6174\ : Span4Mux_v
    port map (
            O => \N__29268\,
            I => \N__29265\
        );

    \I__6173\ : Odrv4
    port map (
            O => \N__29265\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_8\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__29262\,
            I => \N__29258\
        );

    \I__6171\ : InMux
    port map (
            O => \N__29261\,
            I => \N__29254\
        );

    \I__6170\ : InMux
    port map (
            O => \N__29258\,
            I => \N__29249\
        );

    \I__6169\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29249\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__29254\,
            I => \PWMInstance3.periodCounterZ0Z_8\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__29249\,
            I => \PWMInstance3.periodCounterZ0Z_8\
        );

    \I__6166\ : CascadeMux
    port map (
            O => \N__29244\,
            I => \N__29239\
        );

    \I__6165\ : InMux
    port map (
            O => \N__29243\,
            I => \N__29236\
        );

    \I__6164\ : InMux
    port map (
            O => \N__29242\,
            I => \N__29233\
        );

    \I__6163\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29230\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__29236\,
            I => \PWMInstance3.periodCounterZ0Z_9\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__29233\,
            I => \PWMInstance3.periodCounterZ0Z_9\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__29230\,
            I => \PWMInstance3.periodCounterZ0Z_9\
        );

    \I__6159\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29220\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__29220\,
            I => \N__29217\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__29217\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_9\
        );

    \I__6156\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29211\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__29211\,
            I => \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_2\
        );

    \I__6154\ : InMux
    port map (
            O => \N__29208\,
            I => \N__29205\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__29205\,
            I => \N__29202\
        );

    \I__6152\ : Odrv4
    port map (
            O => \N__29202\,
            I => \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_2\
        );

    \I__6151\ : InMux
    port map (
            O => \N__29199\,
            I => \N__29196\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__29196\,
            I => \N__29193\
        );

    \I__6149\ : Span4Mux_v
    port map (
            O => \N__29193\,
            I => \N__29190\
        );

    \I__6148\ : Odrv4
    port map (
            O => \N__29190\,
            I => \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_2\
        );

    \I__6147\ : InMux
    port map (
            O => \N__29187\,
            I => \N__29184\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__29184\,
            I => \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_2\
        );

    \I__6145\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29178\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__29178\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_2\
        );

    \I__6143\ : CascadeMux
    port map (
            O => \N__29175\,
            I => \N__29171\
        );

    \I__6142\ : InMux
    port map (
            O => \N__29174\,
            I => \N__29167\
        );

    \I__6141\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29164\
        );

    \I__6140\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29161\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__29167\,
            I => \PWMInstance3.periodCounterZ0Z_15\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__29164\,
            I => \PWMInstance3.periodCounterZ0Z_15\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__29161\,
            I => \PWMInstance3.periodCounterZ0Z_15\
        );

    \I__6136\ : InMux
    port map (
            O => \N__29154\,
            I => \N__29149\
        );

    \I__6135\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29146\
        );

    \I__6134\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29143\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__29149\,
            I => \N__29140\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__29146\,
            I => \PWMInstance3.periodCounterZ0Z_14\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__29143\,
            I => \PWMInstance3.periodCounterZ0Z_14\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__29140\,
            I => \PWMInstance3.periodCounterZ0Z_14\
        );

    \I__6129\ : InMux
    port map (
            O => \N__29133\,
            I => \N__29130\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__29130\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_14\
        );

    \I__6127\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29124\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__29124\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_15\
        );

    \I__6125\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29118\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__29118\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_13\
        );

    \I__6123\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29112\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__29112\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_12\
        );

    \I__6121\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29104\
        );

    \I__6120\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29101\
        );

    \I__6119\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29098\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__29104\,
            I => \N__29095\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__29101\,
            I => \PWMInstance3.periodCounterZ0Z_12\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__29098\,
            I => \PWMInstance3.periodCounterZ0Z_12\
        );

    \I__6115\ : Odrv4
    port map (
            O => \N__29095\,
            I => \PWMInstance3.periodCounterZ0Z_12\
        );

    \I__6114\ : CascadeMux
    port map (
            O => \N__29088\,
            I => \N__29084\
        );

    \I__6113\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29080\
        );

    \I__6112\ : InMux
    port map (
            O => \N__29084\,
            I => \N__29077\
        );

    \I__6111\ : InMux
    port map (
            O => \N__29083\,
            I => \N__29074\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__29080\,
            I => \PWMInstance3.periodCounterZ0Z_13\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__29077\,
            I => \PWMInstance3.periodCounterZ0Z_13\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__29074\,
            I => \PWMInstance3.periodCounterZ0Z_13\
        );

    \I__6107\ : InMux
    port map (
            O => \N__29067\,
            I => \N__29064\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__29064\,
            I => \N__29061\
        );

    \I__6105\ : Span4Mux_v
    port map (
            O => \N__29061\,
            I => \N__29058\
        );

    \I__6104\ : Odrv4
    port map (
            O => \N__29058\,
            I => \PWMInstance3.un1_periodCounter12_1_0_a2_0_9\
        );

    \I__6103\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29050\
        );

    \I__6102\ : InMux
    port map (
            O => \N__29054\,
            I => \N__29045\
        );

    \I__6101\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29045\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__29050\,
            I => \PWMInstance3.periodCounterZ0Z_0\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__29045\,
            I => \PWMInstance3.periodCounterZ0Z_0\
        );

    \I__6098\ : CascadeMux
    port map (
            O => \N__29040\,
            I => \N__29035\
        );

    \I__6097\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29032\
        );

    \I__6096\ : InMux
    port map (
            O => \N__29038\,
            I => \N__29029\
        );

    \I__6095\ : InMux
    port map (
            O => \N__29035\,
            I => \N__29026\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__29032\,
            I => \PWMInstance3.periodCounterZ0Z_1\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__29029\,
            I => \PWMInstance3.periodCounterZ0Z_1\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__29026\,
            I => \PWMInstance3.periodCounterZ0Z_1\
        );

    \I__6091\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29016\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__29016\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_0\
        );

    \I__6089\ : InMux
    port map (
            O => \N__29013\,
            I => \N__29010\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__29010\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_1\
        );

    \I__6087\ : InMux
    port map (
            O => \N__29007\,
            I => \N__29004\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__29004\,
            I => \N__28999\
        );

    \I__6085\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28996\
        );

    \I__6084\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28993\
        );

    \I__6083\ : Span4Mux_v
    port map (
            O => \N__28999\,
            I => \N__28980\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__28996\,
            I => \N__28980\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__28993\,
            I => \N__28977\
        );

    \I__6080\ : InMux
    port map (
            O => \N__28992\,
            I => \N__28973\
        );

    \I__6079\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28967\
        );

    \I__6078\ : InMux
    port map (
            O => \N__28990\,
            I => \N__28967\
        );

    \I__6077\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28962\
        );

    \I__6076\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28962\
        );

    \I__6075\ : InMux
    port map (
            O => \N__28987\,
            I => \N__28959\
        );

    \I__6074\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28956\
        );

    \I__6073\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28953\
        );

    \I__6072\ : Span4Mux_v
    port map (
            O => \N__28980\,
            I => \N__28947\
        );

    \I__6071\ : Span4Mux_v
    port map (
            O => \N__28977\,
            I => \N__28947\
        );

    \I__6070\ : InMux
    port map (
            O => \N__28976\,
            I => \N__28944\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__28973\,
            I => \N__28940\
        );

    \I__6068\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28937\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__28967\,
            I => \N__28934\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__28962\,
            I => \N__28925\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__28959\,
            I => \N__28925\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__28956\,
            I => \N__28925\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__28953\,
            I => \N__28925\
        );

    \I__6062\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28922\
        );

    \I__6061\ : Span4Mux_h
    port map (
            O => \N__28947\,
            I => \N__28919\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__28944\,
            I => \N__28916\
        );

    \I__6059\ : InMux
    port map (
            O => \N__28943\,
            I => \N__28913\
        );

    \I__6058\ : Span4Mux_v
    port map (
            O => \N__28940\,
            I => \N__28909\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__28937\,
            I => \N__28904\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__28934\,
            I => \N__28904\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__28925\,
            I => \N__28899\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__28922\,
            I => \N__28899\
        );

    \I__6053\ : Span4Mux_h
    port map (
            O => \N__28919\,
            I => \N__28892\
        );

    \I__6052\ : Span4Mux_v
    port map (
            O => \N__28916\,
            I => \N__28892\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28892\
        );

    \I__6050\ : InMux
    port map (
            O => \N__28912\,
            I => \N__28889\
        );

    \I__6049\ : Span4Mux_h
    port map (
            O => \N__28909\,
            I => \N__28882\
        );

    \I__6048\ : Span4Mux_v
    port map (
            O => \N__28904\,
            I => \N__28882\
        );

    \I__6047\ : Span4Mux_v
    port map (
            O => \N__28899\,
            I => \N__28882\
        );

    \I__6046\ : Odrv4
    port map (
            O => \N__28892\,
            I => \dataWriteZ0Z_8\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__28889\,
            I => \dataWriteZ0Z_8\
        );

    \I__6044\ : Odrv4
    port map (
            O => \N__28882\,
            I => \dataWriteZ0Z_8\
        );

    \I__6043\ : InMux
    port map (
            O => \N__28875\,
            I => \N__28867\
        );

    \I__6042\ : CascadeMux
    port map (
            O => \N__28874\,
            I => \N__28863\
        );

    \I__6041\ : InMux
    port map (
            O => \N__28873\,
            I => \N__28858\
        );

    \I__6040\ : InMux
    port map (
            O => \N__28872\,
            I => \N__28855\
        );

    \I__6039\ : InMux
    port map (
            O => \N__28871\,
            I => \N__28851\
        );

    \I__6038\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28848\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28844\
        );

    \I__6036\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28839\
        );

    \I__6035\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28839\
        );

    \I__6034\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28834\
        );

    \I__6033\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28834\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28830\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__28855\,
            I => \N__28827\
        );

    \I__6030\ : InMux
    port map (
            O => \N__28854\,
            I => \N__28824\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__28851\,
            I => \N__28820\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__28848\,
            I => \N__28816\
        );

    \I__6027\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28813\
        );

    \I__6026\ : Span4Mux_v
    port map (
            O => \N__28844\,
            I => \N__28808\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__28839\,
            I => \N__28808\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__28834\,
            I => \N__28805\
        );

    \I__6023\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28802\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__28830\,
            I => \N__28797\
        );

    \I__6021\ : Span4Mux_h
    port map (
            O => \N__28827\,
            I => \N__28794\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__28824\,
            I => \N__28791\
        );

    \I__6019\ : InMux
    port map (
            O => \N__28823\,
            I => \N__28788\
        );

    \I__6018\ : Span4Mux_v
    port map (
            O => \N__28820\,
            I => \N__28785\
        );

    \I__6017\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28782\
        );

    \I__6016\ : Span4Mux_v
    port map (
            O => \N__28816\,
            I => \N__28779\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__28813\,
            I => \N__28776\
        );

    \I__6014\ : Span4Mux_h
    port map (
            O => \N__28808\,
            I => \N__28769\
        );

    \I__6013\ : Span4Mux_h
    port map (
            O => \N__28805\,
            I => \N__28769\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28769\
        );

    \I__6011\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28766\
        );

    \I__6010\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28763\
        );

    \I__6009\ : Span4Mux_h
    port map (
            O => \N__28797\,
            I => \N__28760\
        );

    \I__6008\ : Span4Mux_h
    port map (
            O => \N__28794\,
            I => \N__28753\
        );

    \I__6007\ : Span4Mux_v
    port map (
            O => \N__28791\,
            I => \N__28753\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__28788\,
            I => \N__28753\
        );

    \I__6005\ : Sp12to4
    port map (
            O => \N__28785\,
            I => \N__28748\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__28782\,
            I => \N__28748\
        );

    \I__6003\ : Span4Mux_h
    port map (
            O => \N__28779\,
            I => \N__28737\
        );

    \I__6002\ : Span4Mux_h
    port map (
            O => \N__28776\,
            I => \N__28737\
        );

    \I__6001\ : Span4Mux_h
    port map (
            O => \N__28769\,
            I => \N__28737\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__28766\,
            I => \N__28737\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__28763\,
            I => \N__28737\
        );

    \I__5998\ : Odrv4
    port map (
            O => \N__28760\,
            I => \dataWriteZ0Z_12\
        );

    \I__5997\ : Odrv4
    port map (
            O => \N__28753\,
            I => \dataWriteZ0Z_12\
        );

    \I__5996\ : Odrv12
    port map (
            O => \N__28748\,
            I => \dataWriteZ0Z_12\
        );

    \I__5995\ : Odrv4
    port map (
            O => \N__28737\,
            I => \dataWriteZ0Z_12\
        );

    \I__5994\ : InMux
    port map (
            O => \N__28728\,
            I => \N__28720\
        );

    \I__5993\ : InMux
    port map (
            O => \N__28727\,
            I => \N__28716\
        );

    \I__5992\ : InMux
    port map (
            O => \N__28726\,
            I => \N__28712\
        );

    \I__5991\ : InMux
    port map (
            O => \N__28725\,
            I => \N__28708\
        );

    \I__5990\ : InMux
    port map (
            O => \N__28724\,
            I => \N__28705\
        );

    \I__5989\ : InMux
    port map (
            O => \N__28723\,
            I => \N__28700\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__28720\,
            I => \N__28696\
        );

    \I__5987\ : InMux
    port map (
            O => \N__28719\,
            I => \N__28693\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__28716\,
            I => \N__28690\
        );

    \I__5985\ : InMux
    port map (
            O => \N__28715\,
            I => \N__28687\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__28712\,
            I => \N__28681\
        );

    \I__5983\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28678\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__28708\,
            I => \N__28674\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28671\
        );

    \I__5980\ : InMux
    port map (
            O => \N__28704\,
            I => \N__28668\
        );

    \I__5979\ : InMux
    port map (
            O => \N__28703\,
            I => \N__28665\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__28700\,
            I => \N__28662\
        );

    \I__5977\ : InMux
    port map (
            O => \N__28699\,
            I => \N__28659\
        );

    \I__5976\ : Span4Mux_v
    port map (
            O => \N__28696\,
            I => \N__28654\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__28693\,
            I => \N__28654\
        );

    \I__5974\ : Span4Mux_h
    port map (
            O => \N__28690\,
            I => \N__28649\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__28687\,
            I => \N__28649\
        );

    \I__5972\ : InMux
    port map (
            O => \N__28686\,
            I => \N__28642\
        );

    \I__5971\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28642\
        );

    \I__5970\ : InMux
    port map (
            O => \N__28684\,
            I => \N__28642\
        );

    \I__5969\ : Span4Mux_v
    port map (
            O => \N__28681\,
            I => \N__28639\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__28678\,
            I => \N__28636\
        );

    \I__5967\ : InMux
    port map (
            O => \N__28677\,
            I => \N__28633\
        );

    \I__5966\ : Span4Mux_h
    port map (
            O => \N__28674\,
            I => \N__28630\
        );

    \I__5965\ : Span4Mux_v
    port map (
            O => \N__28671\,
            I => \N__28623\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__28668\,
            I => \N__28623\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__28665\,
            I => \N__28623\
        );

    \I__5962\ : Span4Mux_v
    port map (
            O => \N__28662\,
            I => \N__28620\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__28659\,
            I => \N__28617\
        );

    \I__5960\ : Span4Mux_h
    port map (
            O => \N__28654\,
            I => \N__28610\
        );

    \I__5959\ : Span4Mux_h
    port map (
            O => \N__28649\,
            I => \N__28610\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__28642\,
            I => \N__28610\
        );

    \I__5957\ : Span4Mux_h
    port map (
            O => \N__28639\,
            I => \N__28603\
        );

    \I__5956\ : Span4Mux_v
    port map (
            O => \N__28636\,
            I => \N__28603\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__28633\,
            I => \N__28603\
        );

    \I__5954\ : Span4Mux_h
    port map (
            O => \N__28630\,
            I => \N__28598\
        );

    \I__5953\ : Span4Mux_h
    port map (
            O => \N__28623\,
            I => \N__28598\
        );

    \I__5952\ : Span4Mux_h
    port map (
            O => \N__28620\,
            I => \N__28591\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__28617\,
            I => \N__28591\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__28610\,
            I => \N__28591\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__28603\,
            I => \dataWriteZ0Z_13\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__28598\,
            I => \dataWriteZ0Z_13\
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__28591\,
            I => \dataWriteZ0Z_13\
        );

    \I__5946\ : InMux
    port map (
            O => \N__28584\,
            I => \N__28581\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__28581\,
            I => \N__28573\
        );

    \I__5944\ : InMux
    port map (
            O => \N__28580\,
            I => \N__28569\
        );

    \I__5943\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28566\
        );

    \I__5942\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28560\
        );

    \I__5941\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28560\
        );

    \I__5940\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28554\
        );

    \I__5939\ : Span4Mux_v
    port map (
            O => \N__28573\,
            I => \N__28551\
        );

    \I__5938\ : InMux
    port map (
            O => \N__28572\,
            I => \N__28548\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__28569\,
            I => \N__28545\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__28566\,
            I => \N__28542\
        );

    \I__5935\ : InMux
    port map (
            O => \N__28565\,
            I => \N__28538\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__28560\,
            I => \N__28535\
        );

    \I__5933\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28532\
        );

    \I__5932\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28529\
        );

    \I__5931\ : InMux
    port map (
            O => \N__28557\,
            I => \N__28524\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__28554\,
            I => \N__28520\
        );

    \I__5929\ : Span4Mux_h
    port map (
            O => \N__28551\,
            I => \N__28515\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__28548\,
            I => \N__28515\
        );

    \I__5927\ : Span4Mux_v
    port map (
            O => \N__28545\,
            I => \N__28510\
        );

    \I__5926\ : Span4Mux_v
    port map (
            O => \N__28542\,
            I => \N__28510\
        );

    \I__5925\ : InMux
    port map (
            O => \N__28541\,
            I => \N__28507\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__28538\,
            I => \N__28503\
        );

    \I__5923\ : Span4Mux_h
    port map (
            O => \N__28535\,
            I => \N__28496\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__28532\,
            I => \N__28496\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__28529\,
            I => \N__28496\
        );

    \I__5920\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28491\
        );

    \I__5919\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28491\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28488\
        );

    \I__5917\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28485\
        );

    \I__5916\ : Span4Mux_h
    port map (
            O => \N__28520\,
            I => \N__28482\
        );

    \I__5915\ : Span4Mux_h
    port map (
            O => \N__28515\,
            I => \N__28479\
        );

    \I__5914\ : Span4Mux_h
    port map (
            O => \N__28510\,
            I => \N__28476\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__28507\,
            I => \N__28473\
        );

    \I__5912\ : InMux
    port map (
            O => \N__28506\,
            I => \N__28470\
        );

    \I__5911\ : Span4Mux_v
    port map (
            O => \N__28503\,
            I => \N__28463\
        );

    \I__5910\ : Span4Mux_h
    port map (
            O => \N__28496\,
            I => \N__28463\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__28491\,
            I => \N__28463\
        );

    \I__5908\ : Span4Mux_v
    port map (
            O => \N__28488\,
            I => \N__28458\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__28485\,
            I => \N__28458\
        );

    \I__5906\ : Span4Mux_h
    port map (
            O => \N__28482\,
            I => \N__28453\
        );

    \I__5905\ : Span4Mux_v
    port map (
            O => \N__28479\,
            I => \N__28453\
        );

    \I__5904\ : Span4Mux_h
    port map (
            O => \N__28476\,
            I => \N__28444\
        );

    \I__5903\ : Span4Mux_v
    port map (
            O => \N__28473\,
            I => \N__28444\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__28470\,
            I => \N__28444\
        );

    \I__5901\ : Span4Mux_v
    port map (
            O => \N__28463\,
            I => \N__28444\
        );

    \I__5900\ : Odrv4
    port map (
            O => \N__28458\,
            I => \dataWriteZ0Z_9\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__28453\,
            I => \dataWriteZ0Z_9\
        );

    \I__5898\ : Odrv4
    port map (
            O => \N__28444\,
            I => \dataWriteZ0Z_9\
        );

    \I__5897\ : CascadeMux
    port map (
            O => \N__28437\,
            I => \N__28432\
        );

    \I__5896\ : InMux
    port map (
            O => \N__28436\,
            I => \N__28429\
        );

    \I__5895\ : InMux
    port map (
            O => \N__28435\,
            I => \N__28426\
        );

    \I__5894\ : InMux
    port map (
            O => \N__28432\,
            I => \N__28423\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__28429\,
            I => \PWMInstance3.periodCounterZ0Z_5\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__28426\,
            I => \PWMInstance3.periodCounterZ0Z_5\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__28423\,
            I => \PWMInstance3.periodCounterZ0Z_5\
        );

    \I__5890\ : CascadeMux
    port map (
            O => \N__28416\,
            I => \N__28412\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__28415\,
            I => \N__28408\
        );

    \I__5888\ : InMux
    port map (
            O => \N__28412\,
            I => \N__28405\
        );

    \I__5887\ : InMux
    port map (
            O => \N__28411\,
            I => \N__28402\
        );

    \I__5886\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28399\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__28405\,
            I => \N__28396\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__28402\,
            I => \PWMInstance3.periodCounterZ0Z_11\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__28399\,
            I => \PWMInstance3.periodCounterZ0Z_11\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__28396\,
            I => \PWMInstance3.periodCounterZ0Z_11\
        );

    \I__5881\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28386\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__28386\,
            I => \N__28383\
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__28383\,
            I => \PWMInstance3.un1_periodCounter12_1_0_a2_0_10\
        );

    \I__5878\ : InMux
    port map (
            O => \N__28380\,
            I => \N__28377\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__28377\,
            I => \N__28374\
        );

    \I__5876\ : Span4Mux_h
    port map (
            O => \N__28374\,
            I => \N__28371\
        );

    \I__5875\ : Odrv4
    port map (
            O => \N__28371\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_3\
        );

    \I__5874\ : CascadeMux
    port map (
            O => \N__28368\,
            I => \N__28363\
        );

    \I__5873\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28360\
        );

    \I__5872\ : InMux
    port map (
            O => \N__28366\,
            I => \N__28355\
        );

    \I__5871\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28355\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__28360\,
            I => \PWMInstance3.periodCounterZ0Z_3\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__28355\,
            I => \PWMInstance3.periodCounterZ0Z_3\
        );

    \I__5868\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28345\
        );

    \I__5867\ : InMux
    port map (
            O => \N__28349\,
            I => \N__28342\
        );

    \I__5866\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28339\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__28345\,
            I => \PWMInstance3.periodCounterZ0Z_2\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__28342\,
            I => \PWMInstance3.periodCounterZ0Z_2\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__28339\,
            I => \PWMInstance3.periodCounterZ0Z_2\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__28332\,
            I => \OutReg_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__5861\ : InMux
    port map (
            O => \N__28329\,
            I => \N__28326\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__28326\,
            I => \N__28323\
        );

    \I__5859\ : Span4Mux_v
    port map (
            O => \N__28323\,
            I => \N__28320\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__28320\,
            I => \OutReg_esr_RNO_2Z0Z_6\
        );

    \I__5857\ : CascadeMux
    port map (
            O => \N__28317\,
            I => \OutReg_esr_RNO_0Z0Z_6_cascade_\
        );

    \I__5856\ : InMux
    port map (
            O => \N__28314\,
            I => \N__28311\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__28311\,
            I => \N__28308\
        );

    \I__5854\ : Odrv4
    port map (
            O => \N__28308\,
            I => \OutRegZ0Z_6\
        );

    \I__5853\ : InMux
    port map (
            O => \N__28305\,
            I => \N__28301\
        );

    \I__5852\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28297\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__28301\,
            I => \N__28294\
        );

    \I__5850\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28291\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28288\
        );

    \I__5848\ : Span4Mux_v
    port map (
            O => \N__28294\,
            I => \N__28283\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__28291\,
            I => \N__28283\
        );

    \I__5846\ : Span4Mux_v
    port map (
            O => \N__28288\,
            I => \N__28280\
        );

    \I__5845\ : Span4Mux_v
    port map (
            O => \N__28283\,
            I => \N__28277\
        );

    \I__5844\ : Span4Mux_h
    port map (
            O => \N__28280\,
            I => \N__28274\
        );

    \I__5843\ : Odrv4
    port map (
            O => \N__28277\,
            I => \dataRead2_6\
        );

    \I__5842\ : Odrv4
    port map (
            O => \N__28274\,
            I => \dataRead2_6\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__28269\,
            I => \N__28266\
        );

    \I__5840\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28262\
        );

    \I__5839\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28259\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__28262\,
            I => \N__28255\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__28259\,
            I => \N__28252\
        );

    \I__5836\ : InMux
    port map (
            O => \N__28258\,
            I => \N__28249\
        );

    \I__5835\ : Span4Mux_v
    port map (
            O => \N__28255\,
            I => \N__28246\
        );

    \I__5834\ : Span4Mux_v
    port map (
            O => \N__28252\,
            I => \N__28241\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__28249\,
            I => \N__28241\
        );

    \I__5832\ : Span4Mux_h
    port map (
            O => \N__28246\,
            I => \N__28236\
        );

    \I__5831\ : Span4Mux_h
    port map (
            O => \N__28241\,
            I => \N__28236\
        );

    \I__5830\ : Odrv4
    port map (
            O => \N__28236\,
            I => \dataRead3_6\
        );

    \I__5829\ : InMux
    port map (
            O => \N__28233\,
            I => \N__28230\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__28230\,
            I => \OutReg_0_4_i_m3_ns_1_6\
        );

    \I__5827\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28223\
        );

    \I__5826\ : CascadeMux
    port map (
            O => \N__28226\,
            I => \N__28219\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__28223\,
            I => \N__28216\
        );

    \I__5824\ : CascadeMux
    port map (
            O => \N__28222\,
            I => \N__28213\
        );

    \I__5823\ : InMux
    port map (
            O => \N__28219\,
            I => \N__28210\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__28216\,
            I => \N__28207\
        );

    \I__5821\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28204\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__28210\,
            I => \N__28201\
        );

    \I__5819\ : Span4Mux_h
    port map (
            O => \N__28207\,
            I => \N__28198\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__28204\,
            I => \dataRead5_14\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__28201\,
            I => \dataRead5_14\
        );

    \I__5816\ : Odrv4
    port map (
            O => \N__28198\,
            I => \dataRead5_14\
        );

    \I__5815\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28186\
        );

    \I__5814\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28183\
        );

    \I__5813\ : CascadeMux
    port map (
            O => \N__28189\,
            I => \N__28180\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__28186\,
            I => \N__28177\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__28183\,
            I => \N__28174\
        );

    \I__5810\ : InMux
    port map (
            O => \N__28180\,
            I => \N__28171\
        );

    \I__5809\ : Span4Mux_h
    port map (
            O => \N__28177\,
            I => \N__28168\
        );

    \I__5808\ : Odrv4
    port map (
            O => \N__28174\,
            I => \dataRead1_14\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__28171\,
            I => \dataRead1_14\
        );

    \I__5806\ : Odrv4
    port map (
            O => \N__28168\,
            I => \dataRead1_14\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__28161\,
            I => \OutReg_0_5_i_m3_ns_1_14_cascade_\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__28158\,
            I => \OutReg_esr_RNO_2Z0Z_14_cascade_\
        );

    \I__5803\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28152\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__28152\,
            I => \N__28149\
        );

    \I__5801\ : Odrv12
    port map (
            O => \N__28149\,
            I => \OutReg_esr_RNO_1Z0Z_14\
        );

    \I__5800\ : InMux
    port map (
            O => \N__28146\,
            I => \N__28143\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__28143\,
            I => \OutReg_esr_RNO_0Z0Z_14\
        );

    \I__5798\ : CascadeMux
    port map (
            O => \N__28140\,
            I => \N__28134\
        );

    \I__5797\ : CascadeMux
    port map (
            O => \N__28139\,
            I => \N__28129\
        );

    \I__5796\ : InMux
    port map (
            O => \N__28138\,
            I => \N__28123\
        );

    \I__5795\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28118\
        );

    \I__5794\ : InMux
    port map (
            O => \N__28134\,
            I => \N__28118\
        );

    \I__5793\ : CascadeMux
    port map (
            O => \N__28133\,
            I => \N__28115\
        );

    \I__5792\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28112\
        );

    \I__5791\ : InMux
    port map (
            O => \N__28129\,
            I => \N__28109\
        );

    \I__5790\ : InMux
    port map (
            O => \N__28128\,
            I => \N__28106\
        );

    \I__5789\ : InMux
    port map (
            O => \N__28127\,
            I => \N__28103\
        );

    \I__5788\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28098\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__28123\,
            I => \N__28095\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__28118\,
            I => \N__28092\
        );

    \I__5785\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28089\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__28112\,
            I => \N__28084\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__28109\,
            I => \N__28084\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__28106\,
            I => \N__28081\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__28103\,
            I => \N__28078\
        );

    \I__5780\ : InMux
    port map (
            O => \N__28102\,
            I => \N__28075\
        );

    \I__5779\ : InMux
    port map (
            O => \N__28101\,
            I => \N__28072\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__28098\,
            I => \N__28067\
        );

    \I__5777\ : Span4Mux_v
    port map (
            O => \N__28095\,
            I => \N__28067\
        );

    \I__5776\ : Span4Mux_v
    port map (
            O => \N__28092\,
            I => \N__28062\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__28089\,
            I => \N__28062\
        );

    \I__5774\ : Span12Mux_s7_v
    port map (
            O => \N__28084\,
            I => \N__28059\
        );

    \I__5773\ : Odrv4
    port map (
            O => \N__28081\,
            I => \data_received_2_repZ0Z1\
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__28078\,
            I => \data_received_2_repZ0Z1\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__28075\,
            I => \data_received_2_repZ0Z1\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__28072\,
            I => \data_received_2_repZ0Z1\
        );

    \I__5769\ : Odrv4
    port map (
            O => \N__28067\,
            I => \data_received_2_repZ0Z1\
        );

    \I__5768\ : Odrv4
    port map (
            O => \N__28062\,
            I => \data_received_2_repZ0Z1\
        );

    \I__5767\ : Odrv12
    port map (
            O => \N__28059\,
            I => \data_received_2_repZ0Z1\
        );

    \I__5766\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28039\
        );

    \I__5765\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28036\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__28042\,
            I => \N__28033\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__28039\,
            I => \N__28028\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__28036\,
            I => \N__28028\
        );

    \I__5761\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28025\
        );

    \I__5760\ : Span4Mux_v
    port map (
            O => \N__28028\,
            I => \N__28022\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__28025\,
            I => \dataRead4_3\
        );

    \I__5758\ : Odrv4
    port map (
            O => \N__28022\,
            I => \dataRead4_3\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__28017\,
            I => \N__28009\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__28016\,
            I => \N__28005\
        );

    \I__5755\ : InMux
    port map (
            O => \N__28015\,
            I => \N__28000\
        );

    \I__5754\ : InMux
    port map (
            O => \N__28014\,
            I => \N__28000\
        );

    \I__5753\ : InMux
    port map (
            O => \N__28013\,
            I => \N__27997\
        );

    \I__5752\ : InMux
    port map (
            O => \N__28012\,
            I => \N__27993\
        );

    \I__5751\ : InMux
    port map (
            O => \N__28009\,
            I => \N__27990\
        );

    \I__5750\ : InMux
    port map (
            O => \N__28008\,
            I => \N__27986\
        );

    \I__5749\ : InMux
    port map (
            O => \N__28005\,
            I => \N__27983\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__28000\,
            I => \N__27978\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__27997\,
            I => \N__27978\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__27996\,
            I => \N__27973\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__27993\,
            I => \N__27970\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__27990\,
            I => \N__27967\
        );

    \I__5743\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27964\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__27986\,
            I => \N__27961\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__27983\,
            I => \N__27958\
        );

    \I__5740\ : Span4Mux_v
    port map (
            O => \N__27978\,
            I => \N__27955\
        );

    \I__5739\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27952\
        );

    \I__5738\ : InMux
    port map (
            O => \N__27976\,
            I => \N__27949\
        );

    \I__5737\ : InMux
    port map (
            O => \N__27973\,
            I => \N__27946\
        );

    \I__5736\ : Span4Mux_v
    port map (
            O => \N__27970\,
            I => \N__27941\
        );

    \I__5735\ : Span4Mux_v
    port map (
            O => \N__27967\,
            I => \N__27941\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__27964\,
            I => \N__27936\
        );

    \I__5733\ : Span4Mux_s2_v
    port map (
            O => \N__27961\,
            I => \N__27936\
        );

    \I__5732\ : Span4Mux_v
    port map (
            O => \N__27958\,
            I => \N__27931\
        );

    \I__5731\ : Span4Mux_h
    port map (
            O => \N__27955\,
            I => \N__27931\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__27952\,
            I => \data_received_0_repZ0Z1\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__27949\,
            I => \data_received_0_repZ0Z1\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__27946\,
            I => \data_received_0_repZ0Z1\
        );

    \I__5727\ : Odrv4
    port map (
            O => \N__27941\,
            I => \data_received_0_repZ0Z1\
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__27936\,
            I => \data_received_0_repZ0Z1\
        );

    \I__5725\ : Odrv4
    port map (
            O => \N__27931\,
            I => \data_received_0_repZ0Z1\
        );

    \I__5724\ : InMux
    port map (
            O => \N__27918\,
            I => \N__27914\
        );

    \I__5723\ : InMux
    port map (
            O => \N__27917\,
            I => \N__27910\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__27914\,
            I => \N__27907\
        );

    \I__5721\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27904\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__27910\,
            I => \N__27901\
        );

    \I__5719\ : Span4Mux_h
    port map (
            O => \N__27907\,
            I => \N__27898\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__27904\,
            I => \N__27895\
        );

    \I__5717\ : Span4Mux_v
    port map (
            O => \N__27901\,
            I => \N__27892\
        );

    \I__5716\ : Span4Mux_v
    port map (
            O => \N__27898\,
            I => \N__27889\
        );

    \I__5715\ : Span4Mux_h
    port map (
            O => \N__27895\,
            I => \N__27884\
        );

    \I__5714\ : Span4Mux_h
    port map (
            O => \N__27892\,
            I => \N__27884\
        );

    \I__5713\ : Odrv4
    port map (
            O => \N__27889\,
            I => \dataRead5_3\
        );

    \I__5712\ : Odrv4
    port map (
            O => \N__27884\,
            I => \dataRead5_3\
        );

    \I__5711\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27875\
        );

    \I__5710\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27871\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__27875\,
            I => \N__27868\
        );

    \I__5708\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27865\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__27871\,
            I => \N__27860\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__27868\,
            I => \N__27860\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__27865\,
            I => \N__27857\
        );

    \I__5704\ : Span4Mux_v
    port map (
            O => \N__27860\,
            I => \N__27854\
        );

    \I__5703\ : Span4Mux_h
    port map (
            O => \N__27857\,
            I => \N__27851\
        );

    \I__5702\ : Odrv4
    port map (
            O => \N__27854\,
            I => \dataRead1_3\
        );

    \I__5701\ : Odrv4
    port map (
            O => \N__27851\,
            I => \dataRead1_3\
        );

    \I__5700\ : CascadeMux
    port map (
            O => \N__27846\,
            I => \OutReg_0_5_i_m3_ns_1_3_cascade_\
        );

    \I__5699\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27838\
        );

    \I__5698\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27835\
        );

    \I__5697\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27832\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__27838\,
            I => \N__27829\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__27835\,
            I => \N__27824\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__27832\,
            I => \N__27824\
        );

    \I__5693\ : Span12Mux_s10_h
    port map (
            O => \N__27829\,
            I => \N__27819\
        );

    \I__5692\ : Span12Mux_h
    port map (
            O => \N__27824\,
            I => \N__27819\
        );

    \I__5691\ : Odrv12
    port map (
            O => \N__27819\,
            I => \dataRead7_3\
        );

    \I__5690\ : CascadeMux
    port map (
            O => \N__27816\,
            I => \N__27813\
        );

    \I__5689\ : InMux
    port map (
            O => \N__27813\,
            I => \N__27809\
        );

    \I__5688\ : InMux
    port map (
            O => \N__27812\,
            I => \N__27806\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__27809\,
            I => \N__27803\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__27806\,
            I => \N__27800\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__27803\,
            I => \N__27797\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__27800\,
            I => \N__27793\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__27797\,
            I => \N__27790\
        );

    \I__5682\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27787\
        );

    \I__5681\ : Odrv4
    port map (
            O => \N__27793\,
            I => \dataRead6_3\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__27790\,
            I => \dataRead6_3\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__27787\,
            I => \dataRead6_3\
        );

    \I__5678\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27777\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__27777\,
            I => \N__27774\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__27774\,
            I => \OutReg_0_4_i_m3_ns_1_3\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__27771\,
            I => \OutReg_ess_RNO_1Z0Z_3_cascade_\
        );

    \I__5674\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__27765\,
            I => \OutReg_ess_RNO_2Z0Z_3\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__27762\,
            I => \OutReg_ess_RNO_0Z0Z_3_cascade_\
        );

    \I__5671\ : InMux
    port map (
            O => \N__27759\,
            I => \N__27756\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__27756\,
            I => \OutRegZ0Z_3\
        );

    \I__5669\ : InMux
    port map (
            O => \N__27753\,
            I => \N__27750\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__27750\,
            I => \N__27747\
        );

    \I__5667\ : Span4Mux_v
    port map (
            O => \N__27747\,
            I => \N__27744\
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__27744\,
            I => \OutReg_ess_RNO_0Z0Z_4\
        );

    \I__5665\ : InMux
    port map (
            O => \N__27741\,
            I => \N__27737\
        );

    \I__5664\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27734\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__27737\,
            I => \N__27731\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__27734\,
            I => \N__27728\
        );

    \I__5661\ : Span4Mux_h
    port map (
            O => \N__27731\,
            I => \N__27725\
        );

    \I__5660\ : Span4Mux_v
    port map (
            O => \N__27728\,
            I => \N__27721\
        );

    \I__5659\ : Span4Mux_v
    port map (
            O => \N__27725\,
            I => \N__27718\
        );

    \I__5658\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27715\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__27721\,
            I => \dataRead6_6\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__27718\,
            I => \dataRead6_6\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__27715\,
            I => \dataRead6_6\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__27708\,
            I => \N__27705\
        );

    \I__5653\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27701\
        );

    \I__5652\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27697\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__27701\,
            I => \N__27694\
        );

    \I__5650\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27691\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__27697\,
            I => \N__27688\
        );

    \I__5648\ : Span4Mux_h
    port map (
            O => \N__27694\,
            I => \N__27685\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__27691\,
            I => \N__27682\
        );

    \I__5646\ : Span4Mux_v
    port map (
            O => \N__27688\,
            I => \N__27679\
        );

    \I__5645\ : Span4Mux_v
    port map (
            O => \N__27685\,
            I => \N__27674\
        );

    \I__5644\ : Span4Mux_v
    port map (
            O => \N__27682\,
            I => \N__27674\
        );

    \I__5643\ : Odrv4
    port map (
            O => \N__27679\,
            I => \dataRead7_6\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__27674\,
            I => \dataRead7_6\
        );

    \I__5641\ : InMux
    port map (
            O => \N__27669\,
            I => \N__27666\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__27666\,
            I => \N__27663\
        );

    \I__5639\ : Span4Mux_v
    port map (
            O => \N__27663\,
            I => \N__27660\
        );

    \I__5638\ : Odrv4
    port map (
            O => \N__27660\,
            I => \OutReg_0_5_i_m3_ns_1_7\
        );

    \I__5637\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27654\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__27654\,
            I => \N__27651\
        );

    \I__5635\ : Odrv4
    port map (
            O => \N__27651\,
            I => \QuadInstance4.Quad_RNO_0_4_7\
        );

    \I__5634\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27645\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__27645\,
            I => \N__27641\
        );

    \I__5632\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27637\
        );

    \I__5631\ : Span4Mux_h
    port map (
            O => \N__27641\,
            I => \N__27634\
        );

    \I__5630\ : InMux
    port map (
            O => \N__27640\,
            I => \N__27631\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__27637\,
            I => \dataRead4_7\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__27634\,
            I => \dataRead4_7\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__27631\,
            I => \dataRead4_7\
        );

    \I__5626\ : InMux
    port map (
            O => \N__27624\,
            I => \N__27621\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__27621\,
            I => \N__27618\
        );

    \I__5624\ : Span4Mux_v
    port map (
            O => \N__27618\,
            I => \N__27615\
        );

    \I__5623\ : Odrv4
    port map (
            O => \N__27615\,
            I => \OutReg_0_5_i_m3_ns_1_12\
        );

    \I__5622\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27609\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__27609\,
            I => \N__27606\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__27606\,
            I => \QuadInstance4.Quad_RNO_0_4_12\
        );

    \I__5619\ : CascadeMux
    port map (
            O => \N__27603\,
            I => \N__27600\
        );

    \I__5618\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27596\
        );

    \I__5617\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27592\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__27596\,
            I => \N__27589\
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__27595\,
            I => \N__27586\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__27592\,
            I => \N__27583\
        );

    \I__5613\ : Span4Mux_h
    port map (
            O => \N__27589\,
            I => \N__27580\
        );

    \I__5612\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27577\
        );

    \I__5611\ : Odrv12
    port map (
            O => \N__27583\,
            I => \dataRead4_12\
        );

    \I__5610\ : Odrv4
    port map (
            O => \N__27580\,
            I => \dataRead4_12\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__27577\,
            I => \dataRead4_12\
        );

    \I__5608\ : InMux
    port map (
            O => \N__27570\,
            I => \N__27566\
        );

    \I__5607\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27562\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__27566\,
            I => \N__27559\
        );

    \I__5605\ : InMux
    port map (
            O => \N__27565\,
            I => \N__27556\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__27562\,
            I => \N__27553\
        );

    \I__5603\ : Span4Mux_v
    port map (
            O => \N__27559\,
            I => \N__27548\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__27556\,
            I => \N__27548\
        );

    \I__5601\ : Odrv12
    port map (
            O => \N__27553\,
            I => \dataRead4_13\
        );

    \I__5600\ : Odrv4
    port map (
            O => \N__27548\,
            I => \dataRead4_13\
        );

    \I__5599\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27540\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__27540\,
            I => \N__27537\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__27537\,
            I => \N__27534\
        );

    \I__5596\ : Span4Mux_h
    port map (
            O => \N__27534\,
            I => \N__27531\
        );

    \I__5595\ : Odrv4
    port map (
            O => \N__27531\,
            I => \OutReg_0_5_i_m3_ns_1_13\
        );

    \I__5594\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27524\
        );

    \I__5593\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27521\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__27524\,
            I => \N__27518\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__27521\,
            I => \N__27514\
        );

    \I__5590\ : Span4Mux_v
    port map (
            O => \N__27518\,
            I => \N__27511\
        );

    \I__5589\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27508\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__27514\,
            I => \dataRead4_4\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__27511\,
            I => \dataRead4_4\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__27508\,
            I => \dataRead4_4\
        );

    \I__5585\ : CascadeMux
    port map (
            O => \N__27501\,
            I => \QuadInstance4.un1_count_enable_i_a2_0_1_cascade_\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__27498\,
            I => \N__27495\
        );

    \I__5583\ : InMux
    port map (
            O => \N__27495\,
            I => \N__27492\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__27492\,
            I => \N__27489\
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__27489\,
            I => \QuadInstance4.Quad_RNIJUVR1Z0Z_4\
        );

    \I__5580\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27483\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__27483\,
            I => \N__27480\
        );

    \I__5578\ : Span4Mux_h
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__27477\,
            I => \QuadInstance4.delayedCh_AZ0Z_0\
        );

    \I__5576\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27469\
        );

    \I__5575\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27464\
        );

    \I__5574\ : InMux
    port map (
            O => \N__27472\,
            I => \N__27464\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__27469\,
            I => \QuadInstance4.delayedCh_AZ0Z_1\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__27464\,
            I => \QuadInstance4.delayedCh_AZ0Z_1\
        );

    \I__5571\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27456\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__27456\,
            I => \QuadInstance4.delayedCh_AZ0Z_2\
        );

    \I__5569\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27446\
        );

    \I__5568\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27446\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__27451\,
            I => \N__27436\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__27446\,
            I => \N__27433\
        );

    \I__5565\ : CascadeMux
    port map (
            O => \N__27445\,
            I => \N__27428\
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__27444\,
            I => \N__27424\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__27443\,
            I => \N__27419\
        );

    \I__5562\ : CascadeMux
    port map (
            O => \N__27442\,
            I => \N__27416\
        );

    \I__5561\ : CascadeMux
    port map (
            O => \N__27441\,
            I => \N__27412\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__27440\,
            I => \N__27409\
        );

    \I__5559\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27404\
        );

    \I__5558\ : InMux
    port map (
            O => \N__27436\,
            I => \N__27404\
        );

    \I__5557\ : Span12Mux_v
    port map (
            O => \N__27433\,
            I => \N__27401\
        );

    \I__5556\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27398\
        );

    \I__5555\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27393\
        );

    \I__5554\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27393\
        );

    \I__5553\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27386\
        );

    \I__5552\ : InMux
    port map (
            O => \N__27424\,
            I => \N__27386\
        );

    \I__5551\ : InMux
    port map (
            O => \N__27423\,
            I => \N__27386\
        );

    \I__5550\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27377\
        );

    \I__5549\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27377\
        );

    \I__5548\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27377\
        );

    \I__5547\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27377\
        );

    \I__5546\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27372\
        );

    \I__5545\ : InMux
    port map (
            O => \N__27409\,
            I => \N__27372\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__27404\,
            I => \N__27369\
        );

    \I__5543\ : Odrv12
    port map (
            O => \N__27401\,
            I => \QuadInstance4.count_enable\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__27398\,
            I => \QuadInstance4.count_enable\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__27393\,
            I => \QuadInstance4.count_enable\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__27386\,
            I => \QuadInstance4.count_enable\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__27377\,
            I => \QuadInstance4.count_enable\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__27372\,
            I => \QuadInstance4.count_enable\
        );

    \I__5537\ : Odrv4
    port map (
            O => \N__27369\,
            I => \QuadInstance4.count_enable\
        );

    \I__5536\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27348\
        );

    \I__5535\ : CascadeMux
    port map (
            O => \N__27353\,
            I => \N__27339\
        );

    \I__5534\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27333\
        );

    \I__5533\ : InMux
    port map (
            O => \N__27351\,
            I => \N__27333\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__27348\,
            I => \N__27327\
        );

    \I__5531\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27320\
        );

    \I__5530\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27320\
        );

    \I__5529\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27320\
        );

    \I__5528\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27313\
        );

    \I__5527\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27313\
        );

    \I__5526\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27313\
        );

    \I__5525\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27308\
        );

    \I__5524\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27308\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__27333\,
            I => \N__27305\
        );

    \I__5522\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27298\
        );

    \I__5521\ : InMux
    port map (
            O => \N__27331\,
            I => \N__27298\
        );

    \I__5520\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27298\
        );

    \I__5519\ : Odrv12
    port map (
            O => \N__27327\,
            I => \QuadInstance4.un1_count_enable_i_a2_0_1\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__27320\,
            I => \QuadInstance4.un1_count_enable_i_a2_0_1\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__27313\,
            I => \QuadInstance4.un1_count_enable_i_a2_0_1\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__27308\,
            I => \QuadInstance4.un1_count_enable_i_a2_0_1\
        );

    \I__5515\ : Odrv4
    port map (
            O => \N__27305\,
            I => \QuadInstance4.un1_count_enable_i_a2_0_1\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__27298\,
            I => \QuadInstance4.un1_count_enable_i_a2_0_1\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__27285\,
            I => \N__27282\
        );

    \I__5512\ : InMux
    port map (
            O => \N__27282\,
            I => \N__27279\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__27279\,
            I => \QuadInstance4.Quad_RNIN20S1Z0Z_8\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__27276\,
            I => \N__27273\
        );

    \I__5509\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27270\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__27270\,
            I => \N__27267\
        );

    \I__5507\ : Odrv4
    port map (
            O => \N__27267\,
            I => \QuadInstance4.Quad_RNO_0_4_8\
        );

    \I__5506\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27260\
        );

    \I__5505\ : InMux
    port map (
            O => \N__27263\,
            I => \N__27256\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__27260\,
            I => \N__27253\
        );

    \I__5503\ : CascadeMux
    port map (
            O => \N__27259\,
            I => \N__27250\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__27256\,
            I => \N__27247\
        );

    \I__5501\ : Span4Mux_v
    port map (
            O => \N__27253\,
            I => \N__27244\
        );

    \I__5500\ : InMux
    port map (
            O => \N__27250\,
            I => \N__27241\
        );

    \I__5499\ : Odrv12
    port map (
            O => \N__27247\,
            I => \dataRead4_8\
        );

    \I__5498\ : Odrv4
    port map (
            O => \N__27244\,
            I => \dataRead4_8\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__27241\,
            I => \dataRead4_8\
        );

    \I__5496\ : CascadeMux
    port map (
            O => \N__27234\,
            I => \QuadInstance4.count_enable_cascade_\
        );

    \I__5495\ : CascadeMux
    port map (
            O => \N__27231\,
            I => \N__27228\
        );

    \I__5494\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27225\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__27225\,
            I => \QuadInstance4.Quad_RNIHSVR1Z0Z_2\
        );

    \I__5492\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27217\
        );

    \I__5491\ : InMux
    port map (
            O => \N__27221\,
            I => \N__27214\
        );

    \I__5490\ : InMux
    port map (
            O => \N__27220\,
            I => \N__27211\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__27217\,
            I => \N__27206\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__27214\,
            I => \N__27206\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__27211\,
            I => \N__27203\
        );

    \I__5486\ : Span4Mux_v
    port map (
            O => \N__27206\,
            I => \N__27200\
        );

    \I__5485\ : Odrv4
    port map (
            O => \N__27203\,
            I => \dataRead4_1\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__27200\,
            I => \dataRead4_1\
        );

    \I__5483\ : CascadeMux
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__5482\ : InMux
    port map (
            O => \N__27192\,
            I => \N__27189\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__27189\,
            I => \QuadInstance4.Quad_RNIGRVR1Z0Z_1\
        );

    \I__5480\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__27183\,
            I => \QuadInstance4.Quad_RNO_0_4_2\
        );

    \I__5478\ : CascadeMux
    port map (
            O => \N__27180\,
            I => \N__27175\
        );

    \I__5477\ : InMux
    port map (
            O => \N__27179\,
            I => \N__27172\
        );

    \I__5476\ : InMux
    port map (
            O => \N__27178\,
            I => \N__27169\
        );

    \I__5475\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27166\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__27172\,
            I => \dataRead4_2\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__27169\,
            I => \dataRead4_2\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__27166\,
            I => \dataRead4_2\
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__27159\,
            I => \N__27156\
        );

    \I__5470\ : InMux
    port map (
            O => \N__27156\,
            I => \N__27153\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__27153\,
            I => \QuadInstance4.Quad_RNIITVR1Z0Z_3\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__27150\,
            I => \N__27147\
        );

    \I__5467\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27144\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__27144\,
            I => \QuadInstance4.Quad_RNI39TL1Z0Z_13\
        );

    \I__5465\ : InMux
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__27138\,
            I => \QuadInstance4.Quad_RNI4ATL1Z0Z_14\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__27135\,
            I => \N__27131\
        );

    \I__5462\ : InMux
    port map (
            O => \N__27134\,
            I => \N__27128\
        );

    \I__5461\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27125\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__27128\,
            I => \QuadInstance4.delayedCh_BZ0Z_2\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__27125\,
            I => \QuadInstance4.delayedCh_BZ0Z_2\
        );

    \I__5458\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27117\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__27117\,
            I => \N__27114\
        );

    \I__5456\ : IoSpan4Mux
    port map (
            O => \N__27114\,
            I => \N__27111\
        );

    \I__5455\ : Odrv4
    port map (
            O => \N__27111\,
            I => \ch6_B_c\
        );

    \I__5454\ : InMux
    port map (
            O => \N__27108\,
            I => \N__27105\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__27105\,
            I => \N__27102\
        );

    \I__5452\ : Span4Mux_h
    port map (
            O => \N__27102\,
            I => \N__27099\
        );

    \I__5451\ : Span4Mux_v
    port map (
            O => \N__27099\,
            I => \N__27096\
        );

    \I__5450\ : Span4Mux_v
    port map (
            O => \N__27096\,
            I => \N__27093\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__27093\,
            I => \QuadInstance6.delayedCh_BZ0Z_0\
        );

    \I__5448\ : IoInMux
    port map (
            O => \N__27090\,
            I => \N__27087\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__27087\,
            I => \PWM4_obufLegalizeSB_DFFNet\
        );

    \I__5446\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27081\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__27081\,
            I => \N__27078\
        );

    \I__5444\ : Span4Mux_h
    port map (
            O => \N__27078\,
            I => \N__27075\
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__27075\,
            I => \ch1_B_c\
        );

    \I__5442\ : InMux
    port map (
            O => \N__27072\,
            I => \N__27069\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__27069\,
            I => \N__27066\
        );

    \I__5440\ : Span4Mux_v
    port map (
            O => \N__27066\,
            I => \N__27063\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__27063\,
            I => \QuadInstance1.delayedCh_BZ0Z_0\
        );

    \I__5438\ : InMux
    port map (
            O => \N__27060\,
            I => \N__27057\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__27057\,
            I => \QuadInstance4.Quad_RNO_0_4_5\
        );

    \I__5436\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27049\
        );

    \I__5435\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27046\
        );

    \I__5434\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27043\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__27049\,
            I => \dataRead4_5\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__27046\,
            I => \dataRead4_5\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__27043\,
            I => \dataRead4_5\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__27036\,
            I => \N__27033\
        );

    \I__5429\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27030\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__27030\,
            I => \QuadInstance4.Quad_RNIKVVR1Z0Z_5\
        );

    \I__5427\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27024\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__27024\,
            I => \QuadInstance4.Quad_RNI28TL1Z0Z_12\
        );

    \I__5425\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27018\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__27018\,
            I => \N__27015\
        );

    \I__5423\ : Span12Mux_v
    port map (
            O => \N__27015\,
            I => \N__27012\
        );

    \I__5422\ : Odrv12
    port map (
            O => \N__27012\,
            I => \PWMInstance4.un1_periodCounter12_1_0_a2_0\
        );

    \I__5421\ : InMux
    port map (
            O => \N__27009\,
            I => \N__27004\
        );

    \I__5420\ : InMux
    port map (
            O => \N__27008\,
            I => \N__26999\
        );

    \I__5419\ : InMux
    port map (
            O => \N__27007\,
            I => \N__26999\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__27004\,
            I => \PWMInstance4.periodCounterZ0Z_16\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__26999\,
            I => \PWMInstance4.periodCounterZ0Z_16\
        );

    \I__5416\ : InMux
    port map (
            O => \N__26994\,
            I => \N__26989\
        );

    \I__5415\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26986\
        );

    \I__5414\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26983\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__26989\,
            I => \PWMInstance4.periodCounterZ0Z_7\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__26986\,
            I => \PWMInstance4.periodCounterZ0Z_7\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__26983\,
            I => \PWMInstance4.periodCounterZ0Z_7\
        );

    \I__5410\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26967\
        );

    \I__5409\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26967\
        );

    \I__5408\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26967\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__26967\,
            I => \N__26964\
        );

    \I__5406\ : Span12Mux_s9_v
    port map (
            O => \N__26964\,
            I => \N__26961\
        );

    \I__5405\ : Odrv12
    port map (
            O => \N__26961\,
            I => \pwmWriteZ0Z_4\
        );

    \I__5404\ : CEMux
    port map (
            O => \N__26958\,
            I => \N__26955\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__26955\,
            I => \N__26949\
        );

    \I__5402\ : CEMux
    port map (
            O => \N__26954\,
            I => \N__26946\
        );

    \I__5401\ : CEMux
    port map (
            O => \N__26953\,
            I => \N__26943\
        );

    \I__5400\ : CEMux
    port map (
            O => \N__26952\,
            I => \N__26940\
        );

    \I__5399\ : Span4Mux_h
    port map (
            O => \N__26949\,
            I => \N__26935\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__26946\,
            I => \N__26935\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__26943\,
            I => \N__26931\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__26940\,
            I => \N__26928\
        );

    \I__5395\ : Span4Mux_v
    port map (
            O => \N__26935\,
            I => \N__26925\
        );

    \I__5394\ : CEMux
    port map (
            O => \N__26934\,
            I => \N__26922\
        );

    \I__5393\ : Span4Mux_h
    port map (
            O => \N__26931\,
            I => \N__26919\
        );

    \I__5392\ : Span4Mux_h
    port map (
            O => \N__26928\,
            I => \N__26916\
        );

    \I__5391\ : Sp12to4
    port map (
            O => \N__26925\,
            I => \N__26911\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__26922\,
            I => \N__26911\
        );

    \I__5389\ : Odrv4
    port map (
            O => \N__26919\,
            I => \PWMInstance4.pwmWrite_0_4\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__26916\,
            I => \PWMInstance4.pwmWrite_0_4\
        );

    \I__5387\ : Odrv12
    port map (
            O => \N__26911\,
            I => \PWMInstance4.pwmWrite_0_4\
        );

    \I__5386\ : InMux
    port map (
            O => \N__26904\,
            I => \N__26898\
        );

    \I__5385\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26898\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__5383\ : Span12Mux_s10_v
    port map (
            O => \N__26895\,
            I => \N__26892\
        );

    \I__5382\ : Odrv12
    port map (
            O => \N__26892\,
            I => \pwmWrite_fastZ0Z_4\
        );

    \I__5381\ : CascadeMux
    port map (
            O => \N__26889\,
            I => \N__26884\
        );

    \I__5380\ : InMux
    port map (
            O => \N__26888\,
            I => \N__26874\
        );

    \I__5379\ : InMux
    port map (
            O => \N__26887\,
            I => \N__26874\
        );

    \I__5378\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26874\
        );

    \I__5377\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26874\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__26874\,
            I => \PWMInstance4.clkCountZ0Z_1\
        );

    \I__5375\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26859\
        );

    \I__5374\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26859\
        );

    \I__5373\ : InMux
    port map (
            O => \N__26869\,
            I => \N__26859\
        );

    \I__5372\ : InMux
    port map (
            O => \N__26868\,
            I => \N__26859\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__26859\,
            I => \PWMInstance4.clkCountZ0Z_0\
        );

    \I__5370\ : CascadeMux
    port map (
            O => \N__26856\,
            I => \N__26852\
        );

    \I__5369\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26849\
        );

    \I__5368\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26846\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__26849\,
            I => \PWMInstance4.periodCounter12\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__26846\,
            I => \PWMInstance4.periodCounter12\
        );

    \I__5365\ : CascadeMux
    port map (
            O => \N__26841\,
            I => \N__26838\
        );

    \I__5364\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__26835\,
            I => \N__26830\
        );

    \I__5362\ : InMux
    port map (
            O => \N__26834\,
            I => \N__26827\
        );

    \I__5361\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26824\
        );

    \I__5360\ : Span4Mux_v
    port map (
            O => \N__26830\,
            I => \N__26821\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__26827\,
            I => \PWMInstance4.periodCounterZ0Z_15\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__26824\,
            I => \PWMInstance4.periodCounterZ0Z_15\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__26821\,
            I => \PWMInstance4.periodCounterZ0Z_15\
        );

    \I__5356\ : CascadeMux
    port map (
            O => \N__26814\,
            I => \N__26809\
        );

    \I__5355\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26806\
        );

    \I__5354\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26803\
        );

    \I__5353\ : InMux
    port map (
            O => \N__26809\,
            I => \N__26800\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__26806\,
            I => \PWMInstance4.periodCounterZ0Z_1\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__26803\,
            I => \PWMInstance4.periodCounterZ0Z_1\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__26800\,
            I => \PWMInstance4.periodCounterZ0Z_1\
        );

    \I__5349\ : CascadeMux
    port map (
            O => \N__26793\,
            I => \PWMInstance4.periodCounter12_cascade_\
        );

    \I__5348\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__26787\,
            I => \PWMInstance4.un1_periodCounter12_1_0_a2_0_6\
        );

    \I__5346\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26781\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__26781\,
            I => \N__26778\
        );

    \I__5344\ : Odrv4
    port map (
            O => \N__26778\,
            I => \PWMInstance4.un1_periodCounter12_1_0_a2_0_10\
        );

    \I__5343\ : InMux
    port map (
            O => \N__26775\,
            I => \N__26772\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__26772\,
            I => \PWMInstance4.un1_periodCounter12_1_0_a2_0_9\
        );

    \I__5341\ : CascadeMux
    port map (
            O => \N__26769\,
            I => \PWMInstance4.un1_periodCounter12_1_0_a2_0_14_cascade_\
        );

    \I__5340\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26763\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__26763\,
            I => \N__26760\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__26760\,
            I => \PWMInstance4.un1_periodCounter12_1_0_a2_0_12\
        );

    \I__5337\ : CascadeMux
    port map (
            O => \N__26757\,
            I => \N__26754\
        );

    \I__5336\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__26751\,
            I => \N__26743\
        );

    \I__5334\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26740\
        );

    \I__5333\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26737\
        );

    \I__5332\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26732\
        );

    \I__5331\ : InMux
    port map (
            O => \N__26747\,
            I => \N__26732\
        );

    \I__5330\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26729\
        );

    \I__5329\ : Span12Mux_s11_v
    port map (
            O => \N__26743\,
            I => \N__26726\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__26740\,
            I => \PWMInstance4.out_0_sqmuxa\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__26737\,
            I => \PWMInstance4.out_0_sqmuxa\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__26732\,
            I => \PWMInstance4.out_0_sqmuxa\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__26729\,
            I => \PWMInstance4.out_0_sqmuxa\
        );

    \I__5324\ : Odrv12
    port map (
            O => \N__26726\,
            I => \PWMInstance4.out_0_sqmuxa\
        );

    \I__5323\ : InMux
    port map (
            O => \N__26715\,
            I => \PWMInstance3.un1_periodCounter_2_cry_14\
        );

    \I__5322\ : InMux
    port map (
            O => \N__26712\,
            I => \bfn_15_15_0_\
        );

    \I__5321\ : CascadeMux
    port map (
            O => \N__26709\,
            I => \N__26706\
        );

    \I__5320\ : InMux
    port map (
            O => \N__26706\,
            I => \N__26699\
        );

    \I__5319\ : InMux
    port map (
            O => \N__26705\,
            I => \N__26699\
        );

    \I__5318\ : InMux
    port map (
            O => \N__26704\,
            I => \N__26696\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26693\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__26696\,
            I => \PWMInstance3.periodCounterZ0Z_16\
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__26693\,
            I => \PWMInstance3.periodCounterZ0Z_16\
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__26688\,
            I => \N__26685\
        );

    \I__5313\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26680\
        );

    \I__5312\ : InMux
    port map (
            O => \N__26684\,
            I => \N__26677\
        );

    \I__5311\ : InMux
    port map (
            O => \N__26683\,
            I => \N__26674\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__26680\,
            I => \N__26669\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__26677\,
            I => \N__26669\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__26674\,
            I => \PWMInstance4.periodCounterZ0Z_13\
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__26669\,
            I => \PWMInstance4.periodCounterZ0Z_13\
        );

    \I__5306\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26659\
        );

    \I__5305\ : InMux
    port map (
            O => \N__26663\,
            I => \N__26654\
        );

    \I__5304\ : InMux
    port map (
            O => \N__26662\,
            I => \N__26654\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__26659\,
            I => \PWMInstance4.periodCounterZ0Z_0\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__26654\,
            I => \PWMInstance4.periodCounterZ0Z_0\
        );

    \I__5301\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26646\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__26646\,
            I => \N__26643\
        );

    \I__5299\ : Span4Mux_v
    port map (
            O => \N__26643\,
            I => \N__26640\
        );

    \I__5298\ : Odrv4
    port map (
            O => \N__26640\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_0\
        );

    \I__5297\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26634\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__26634\,
            I => \N__26631\
        );

    \I__5295\ : Span12Mux_s4_v
    port map (
            O => \N__26631\,
            I => \N__26628\
        );

    \I__5294\ : Odrv12
    port map (
            O => \N__26628\,
            I => \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_3\
        );

    \I__5293\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26622\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__26622\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_1\
        );

    \I__5291\ : InMux
    port map (
            O => \N__26619\,
            I => \N__26614\
        );

    \I__5290\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26609\
        );

    \I__5289\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26609\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__26614\,
            I => \PWMInstance4.periodCounterZ0Z_6\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__26609\,
            I => \PWMInstance4.periodCounterZ0Z_6\
        );

    \I__5286\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26601\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__26601\,
            I => \N__26598\
        );

    \I__5284\ : Span12Mux_s7_v
    port map (
            O => \N__26598\,
            I => \N__26595\
        );

    \I__5283\ : Odrv12
    port map (
            O => \N__26595\,
            I => \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_3\
        );

    \I__5282\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26589\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__26589\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_6\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__26586\,
            I => \N__26583\
        );

    \I__5279\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26580\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__26580\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_7\
        );

    \I__5277\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__26574\,
            I => \N__26571\
        );

    \I__5275\ : Odrv4
    port map (
            O => \N__26571\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_9\
        );

    \I__5274\ : CascadeMux
    port map (
            O => \N__26568\,
            I => \N__26564\
        );

    \I__5273\ : InMux
    port map (
            O => \N__26567\,
            I => \N__26560\
        );

    \I__5272\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26555\
        );

    \I__5271\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26555\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__26560\,
            I => \PWMInstance4.periodCounterZ0Z_8\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__26555\,
            I => \PWMInstance4.periodCounterZ0Z_8\
        );

    \I__5268\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26545\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__26549\,
            I => \N__26542\
        );

    \I__5266\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26539\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__26545\,
            I => \N__26536\
        );

    \I__5264\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26533\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__26539\,
            I => \PWMInstance4.periodCounterZ0Z_9\
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__26536\,
            I => \PWMInstance4.periodCounterZ0Z_9\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__26533\,
            I => \PWMInstance4.periodCounterZ0Z_9\
        );

    \I__5260\ : InMux
    port map (
            O => \N__26526\,
            I => \N__26523\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__26523\,
            I => \N__26520\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__26520\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_8\
        );

    \I__5257\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26514\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__26514\,
            I => \N__26511\
        );

    \I__5255\ : Span12Mux_s10_v
    port map (
            O => \N__26511\,
            I => \N__26508\
        );

    \I__5254\ : Odrv12
    port map (
            O => \N__26508\,
            I => \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_3\
        );

    \I__5253\ : InMux
    port map (
            O => \N__26505\,
            I => \PWMInstance3.un1_periodCounter_2_cry_5\
        );

    \I__5252\ : InMux
    port map (
            O => \N__26502\,
            I => \PWMInstance3.un1_periodCounter_2_cry_6\
        );

    \I__5251\ : InMux
    port map (
            O => \N__26499\,
            I => \bfn_15_14_0_\
        );

    \I__5250\ : InMux
    port map (
            O => \N__26496\,
            I => \PWMInstance3.un1_periodCounter_2_cry_8\
        );

    \I__5249\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26486\
        );

    \I__5248\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26486\
        );

    \I__5247\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26483\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26480\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__26483\,
            I => \PWMInstance3.periodCounterZ0Z_10\
        );

    \I__5244\ : Odrv4
    port map (
            O => \N__26480\,
            I => \PWMInstance3.periodCounterZ0Z_10\
        );

    \I__5243\ : InMux
    port map (
            O => \N__26475\,
            I => \PWMInstance3.un1_periodCounter_2_cry_9\
        );

    \I__5242\ : InMux
    port map (
            O => \N__26472\,
            I => \PWMInstance3.un1_periodCounter_2_cry_10\
        );

    \I__5241\ : InMux
    port map (
            O => \N__26469\,
            I => \PWMInstance3.un1_periodCounter_2_cry_11\
        );

    \I__5240\ : InMux
    port map (
            O => \N__26466\,
            I => \PWMInstance3.un1_periodCounter_2_cry_12\
        );

    \I__5239\ : InMux
    port map (
            O => \N__26463\,
            I => \PWMInstance3.un1_periodCounter_2_cry_13\
        );

    \I__5238\ : CascadeMux
    port map (
            O => \N__26460\,
            I => \PWMInstance3.un1_periodCounter12_1_0_a2_0_0_cascade_\
        );

    \I__5237\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26454\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__26454\,
            I => \PWMInstance3.un1_periodCounter12_1_0_a2_0_12\
        );

    \I__5235\ : InMux
    port map (
            O => \N__26451\,
            I => \N__26448\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__26448\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_4\
        );

    \I__5233\ : InMux
    port map (
            O => \N__26445\,
            I => \N__26442\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__26442\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_11\
        );

    \I__5231\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26436\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__26436\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_10\
        );

    \I__5229\ : CascadeMux
    port map (
            O => \N__26433\,
            I => \N__26429\
        );

    \I__5228\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26425\
        );

    \I__5227\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26422\
        );

    \I__5226\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26419\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__26425\,
            I => \PWMInstance3.periodCounter12\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__26422\,
            I => \PWMInstance3.periodCounter12\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__26419\,
            I => \PWMInstance3.periodCounter12\
        );

    \I__5222\ : InMux
    port map (
            O => \N__26412\,
            I => \PWMInstance3.un1_periodCounter_2_cry_0\
        );

    \I__5221\ : InMux
    port map (
            O => \N__26409\,
            I => \PWMInstance3.un1_periodCounter_2_cry_1\
        );

    \I__5220\ : InMux
    port map (
            O => \N__26406\,
            I => \PWMInstance3.un1_periodCounter_2_cry_2\
        );

    \I__5219\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26398\
        );

    \I__5218\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26393\
        );

    \I__5217\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26393\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__26398\,
            I => \PWMInstance3.periodCounterZ0Z_4\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__26393\,
            I => \PWMInstance3.periodCounterZ0Z_4\
        );

    \I__5214\ : InMux
    port map (
            O => \N__26388\,
            I => \PWMInstance3.un1_periodCounter_2_cry_3\
        );

    \I__5213\ : InMux
    port map (
            O => \N__26385\,
            I => \PWMInstance3.un1_periodCounter_2_cry_4\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__26382\,
            I => \OutReg_ess_RNO_2Z0Z_7_cascade_\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__26379\,
            I => \OutReg_ess_RNO_0Z0Z_7_cascade_\
        );

    \I__5210\ : InMux
    port map (
            O => \N__26376\,
            I => \N__26371\
        );

    \I__5209\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26368\
        );

    \I__5208\ : InMux
    port map (
            O => \N__26374\,
            I => \N__26365\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__26371\,
            I => \N__26362\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__26368\,
            I => \N__26359\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__26365\,
            I => \N__26356\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__26362\,
            I => \N__26353\
        );

    \I__5203\ : Span4Mux_h
    port map (
            O => \N__26359\,
            I => \N__26350\
        );

    \I__5202\ : Span4Mux_h
    port map (
            O => \N__26356\,
            I => \N__26345\
        );

    \I__5201\ : Span4Mux_v
    port map (
            O => \N__26353\,
            I => \N__26345\
        );

    \I__5200\ : Odrv4
    port map (
            O => \N__26350\,
            I => \dataRead2_7\
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__26345\,
            I => \dataRead2_7\
        );

    \I__5198\ : CascadeMux
    port map (
            O => \N__26340\,
            I => \N__26337\
        );

    \I__5197\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26333\
        );

    \I__5196\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26330\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__26333\,
            I => \N__26326\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__26330\,
            I => \N__26323\
        );

    \I__5193\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26320\
        );

    \I__5192\ : Span4Mux_h
    port map (
            O => \N__26326\,
            I => \N__26317\
        );

    \I__5191\ : Span4Mux_v
    port map (
            O => \N__26323\,
            I => \N__26312\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__26320\,
            I => \N__26312\
        );

    \I__5189\ : Span4Mux_v
    port map (
            O => \N__26317\,
            I => \N__26309\
        );

    \I__5188\ : Odrv4
    port map (
            O => \N__26312\,
            I => \dataRead3_7\
        );

    \I__5187\ : Odrv4
    port map (
            O => \N__26309\,
            I => \dataRead3_7\
        );

    \I__5186\ : InMux
    port map (
            O => \N__26304\,
            I => \N__26300\
        );

    \I__5185\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26297\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__26300\,
            I => \N__26294\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__26297\,
            I => \N__26291\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__26294\,
            I => \N__26288\
        );

    \I__5181\ : Span12Mux_v
    port map (
            O => \N__26291\,
            I => \N__26284\
        );

    \I__5180\ : Span4Mux_v
    port map (
            O => \N__26288\,
            I => \N__26281\
        );

    \I__5179\ : InMux
    port map (
            O => \N__26287\,
            I => \N__26278\
        );

    \I__5178\ : Odrv12
    port map (
            O => \N__26284\,
            I => \dataRead6_7\
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__26281\,
            I => \dataRead6_7\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__26278\,
            I => \dataRead6_7\
        );

    \I__5175\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26267\
        );

    \I__5174\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26264\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__26267\,
            I => \N__26261\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__26264\,
            I => \N__26258\
        );

    \I__5171\ : Span4Mux_v
    port map (
            O => \N__26261\,
            I => \N__26252\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__26258\,
            I => \N__26252\
        );

    \I__5169\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26249\
        );

    \I__5168\ : Span4Mux_h
    port map (
            O => \N__26252\,
            I => \N__26244\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__26249\,
            I => \N__26244\
        );

    \I__5166\ : Span4Mux_v
    port map (
            O => \N__26244\,
            I => \N__26241\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__26241\,
            I => \dataRead7_7\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__26238\,
            I => \OutReg_0_4_i_m3_ns_1_7_cascade_\
        );

    \I__5163\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26232\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__26232\,
            I => \OutReg_ess_RNO_1Z0Z_7\
        );

    \I__5161\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26226\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__26226\,
            I => \N__26223\
        );

    \I__5159\ : Odrv4
    port map (
            O => \N__26223\,
            I => \OutReg_ess_RNO_0Z0Z_9\
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__26220\,
            I => \N__26217\
        );

    \I__5157\ : InMux
    port map (
            O => \N__26217\,
            I => \N__26214\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__26214\,
            I => \N__26211\
        );

    \I__5155\ : Span4Mux_v
    port map (
            O => \N__26211\,
            I => \N__26208\
        );

    \I__5154\ : Odrv4
    port map (
            O => \N__26208\,
            I => \OutRegZ0Z_13\
        );

    \I__5153\ : CascadeMux
    port map (
            O => \N__26205\,
            I => \N__26202\
        );

    \I__5152\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26199\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__26199\,
            I => \N__26196\
        );

    \I__5150\ : Span4Mux_h
    port map (
            O => \N__26196\,
            I => \N__26193\
        );

    \I__5149\ : Odrv4
    port map (
            O => \N__26193\,
            I => \OutRegZ0Z_14\
        );

    \I__5148\ : InMux
    port map (
            O => \N__26190\,
            I => \N__26187\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__26187\,
            I => \PWMInstance3.PWMPulseWidthCountZ0Z_5\
        );

    \I__5146\ : CEMux
    port map (
            O => \N__26184\,
            I => \N__26163\
        );

    \I__5145\ : CEMux
    port map (
            O => \N__26183\,
            I => \N__26163\
        );

    \I__5144\ : CEMux
    port map (
            O => \N__26182\,
            I => \N__26163\
        );

    \I__5143\ : CEMux
    port map (
            O => \N__26181\,
            I => \N__26163\
        );

    \I__5142\ : CEMux
    port map (
            O => \N__26180\,
            I => \N__26163\
        );

    \I__5141\ : CEMux
    port map (
            O => \N__26179\,
            I => \N__26163\
        );

    \I__5140\ : CEMux
    port map (
            O => \N__26178\,
            I => \N__26163\
        );

    \I__5139\ : GlobalMux
    port map (
            O => \N__26163\,
            I => \N__26160\
        );

    \I__5138\ : gio2CtrlBuf
    port map (
            O => \N__26160\,
            I => \N_45_0_g\
        );

    \I__5137\ : SRMux
    port map (
            O => \N__26157\,
            I => \N__26136\
        );

    \I__5136\ : SRMux
    port map (
            O => \N__26156\,
            I => \N__26136\
        );

    \I__5135\ : SRMux
    port map (
            O => \N__26155\,
            I => \N__26136\
        );

    \I__5134\ : SRMux
    port map (
            O => \N__26154\,
            I => \N__26136\
        );

    \I__5133\ : SRMux
    port map (
            O => \N__26153\,
            I => \N__26136\
        );

    \I__5132\ : SRMux
    port map (
            O => \N__26152\,
            I => \N__26136\
        );

    \I__5131\ : SRMux
    port map (
            O => \N__26151\,
            I => \N__26136\
        );

    \I__5130\ : GlobalMux
    port map (
            O => \N__26136\,
            I => \N__26133\
        );

    \I__5129\ : gio2CtrlBuf
    port map (
            O => \N__26133\,
            I => \N_1187_g\
        );

    \I__5128\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26127\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__26127\,
            I => \N__26124\
        );

    \I__5126\ : Odrv12
    port map (
            O => \N__26124\,
            I => \QuadInstance4.Quad_RNO_0_4_13\
        );

    \I__5125\ : InMux
    port map (
            O => \N__26121\,
            I => \N__26118\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__26118\,
            I => \N__26115\
        );

    \I__5123\ : Odrv12
    port map (
            O => \N__26115\,
            I => \QuadInstance7.Quad_RNO_0_7_13\
        );

    \I__5122\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26109\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__26109\,
            I => \N__26104\
        );

    \I__5120\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26101\
        );

    \I__5119\ : CascadeMux
    port map (
            O => \N__26107\,
            I => \N__26098\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__26104\,
            I => \N__26093\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__26101\,
            I => \N__26093\
        );

    \I__5116\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26090\
        );

    \I__5115\ : Span4Mux_h
    port map (
            O => \N__26093\,
            I => \N__26087\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__26090\,
            I => \N__26084\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__26087\,
            I => \dataRead7_13\
        );

    \I__5112\ : Odrv12
    port map (
            O => \N__26084\,
            I => \dataRead7_13\
        );

    \I__5111\ : InMux
    port map (
            O => \N__26079\,
            I => \N__26076\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__26076\,
            I => \N__26073\
        );

    \I__5109\ : Odrv12
    port map (
            O => \N__26073\,
            I => \QuadInstance4.Quad_RNO_0_4_3\
        );

    \I__5108\ : InMux
    port map (
            O => \N__26070\,
            I => \N__26067\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__26067\,
            I => \N__26064\
        );

    \I__5106\ : Span4Mux_h
    port map (
            O => \N__26064\,
            I => \N__26061\
        );

    \I__5105\ : Span4Mux_h
    port map (
            O => \N__26061\,
            I => \N__26058\
        );

    \I__5104\ : Odrv4
    port map (
            O => \N__26058\,
            I => \QuadInstance7.Quad_RNO_0_7_3\
        );

    \I__5103\ : InMux
    port map (
            O => \N__26055\,
            I => \N__26047\
        );

    \I__5102\ : InMux
    port map (
            O => \N__26054\,
            I => \N__26047\
        );

    \I__5101\ : InMux
    port map (
            O => \N__26053\,
            I => \N__26044\
        );

    \I__5100\ : InMux
    port map (
            O => \N__26052\,
            I => \N__26034\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__26047\,
            I => \N__26031\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__26044\,
            I => \N__26028\
        );

    \I__5097\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26025\
        );

    \I__5096\ : CascadeMux
    port map (
            O => \N__26042\,
            I => \N__26022\
        );

    \I__5095\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26015\
        );

    \I__5094\ : InMux
    port map (
            O => \N__26040\,
            I => \N__26015\
        );

    \I__5093\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26015\
        );

    \I__5092\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26008\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__26037\,
            I => \N__26005\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__26034\,
            I => \N__26001\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__26031\,
            I => \N__25994\
        );

    \I__5088\ : Span4Mux_v
    port map (
            O => \N__26028\,
            I => \N__25994\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__26025\,
            I => \N__25994\
        );

    \I__5086\ : InMux
    port map (
            O => \N__26022\,
            I => \N__25991\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__26015\,
            I => \N__25988\
        );

    \I__5084\ : InMux
    port map (
            O => \N__26014\,
            I => \N__25983\
        );

    \I__5083\ : InMux
    port map (
            O => \N__26013\,
            I => \N__25983\
        );

    \I__5082\ : InMux
    port map (
            O => \N__26012\,
            I => \N__25980\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__26011\,
            I => \N__25977\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__26008\,
            I => \N__25966\
        );

    \I__5079\ : InMux
    port map (
            O => \N__26005\,
            I => \N__25961\
        );

    \I__5078\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25961\
        );

    \I__5077\ : Span4Mux_v
    port map (
            O => \N__26001\,
            I => \N__25956\
        );

    \I__5076\ : Span4Mux_h
    port map (
            O => \N__25994\,
            I => \N__25956\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25951\
        );

    \I__5074\ : Span4Mux_v
    port map (
            O => \N__25988\,
            I => \N__25951\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__25983\,
            I => \N__25946\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__25980\,
            I => \N__25946\
        );

    \I__5071\ : InMux
    port map (
            O => \N__25977\,
            I => \N__25943\
        );

    \I__5070\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25936\
        );

    \I__5069\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25936\
        );

    \I__5068\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25936\
        );

    \I__5067\ : CascadeMux
    port map (
            O => \N__25973\,
            I => \N__25932\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__25972\,
            I => \N__25929\
        );

    \I__5065\ : CascadeMux
    port map (
            O => \N__25971\,
            I => \N__25924\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__25970\,
            I => \N__25921\
        );

    \I__5063\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25914\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__25966\,
            I => \N__25907\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__25961\,
            I => \N__25907\
        );

    \I__5060\ : Span4Mux_h
    port map (
            O => \N__25956\,
            I => \N__25907\
        );

    \I__5059\ : Span4Mux_h
    port map (
            O => \N__25951\,
            I => \N__25902\
        );

    \I__5058\ : Span4Mux_v
    port map (
            O => \N__25946\,
            I => \N__25902\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__25943\,
            I => \N__25897\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__25936\,
            I => \N__25897\
        );

    \I__5055\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25888\
        );

    \I__5054\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25888\
        );

    \I__5053\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25888\
        );

    \I__5052\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25888\
        );

    \I__5051\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25877\
        );

    \I__5050\ : InMux
    port map (
            O => \N__25924\,
            I => \N__25877\
        );

    \I__5049\ : InMux
    port map (
            O => \N__25921\,
            I => \N__25877\
        );

    \I__5048\ : InMux
    port map (
            O => \N__25920\,
            I => \N__25877\
        );

    \I__5047\ : InMux
    port map (
            O => \N__25919\,
            I => \N__25877\
        );

    \I__5046\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25872\
        );

    \I__5045\ : InMux
    port map (
            O => \N__25917\,
            I => \N__25872\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__25914\,
            I => \quadWriteZ0Z_7\
        );

    \I__5043\ : Odrv4
    port map (
            O => \N__25907\,
            I => \quadWriteZ0Z_7\
        );

    \I__5042\ : Odrv4
    port map (
            O => \N__25902\,
            I => \quadWriteZ0Z_7\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__25897\,
            I => \quadWriteZ0Z_7\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__25888\,
            I => \quadWriteZ0Z_7\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__25877\,
            I => \quadWriteZ0Z_7\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__25872\,
            I => \quadWriteZ0Z_7\
        );

    \I__5037\ : InMux
    port map (
            O => \N__25857\,
            I => \N__25854\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__25854\,
            I => \N__25851\
        );

    \I__5035\ : Span4Mux_h
    port map (
            O => \N__25851\,
            I => \N__25848\
        );

    \I__5034\ : Span4Mux_h
    port map (
            O => \N__25848\,
            I => \N__25845\
        );

    \I__5033\ : Odrv4
    port map (
            O => \N__25845\,
            I => \QuadInstance7.Quad_RNO_0_6_1\
        );

    \I__5032\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25838\
        );

    \I__5031\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25835\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__25838\,
            I => \N__25831\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__25835\,
            I => \N__25828\
        );

    \I__5028\ : InMux
    port map (
            O => \N__25834\,
            I => \N__25825\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__25831\,
            I => \N__25822\
        );

    \I__5026\ : Sp12to4
    port map (
            O => \N__25828\,
            I => \N__25819\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__25825\,
            I => \N__25816\
        );

    \I__5024\ : Span4Mux_h
    port map (
            O => \N__25822\,
            I => \N__25813\
        );

    \I__5023\ : Odrv12
    port map (
            O => \N__25819\,
            I => \dataRead7_1\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__25816\,
            I => \dataRead7_1\
        );

    \I__5021\ : Odrv4
    port map (
            O => \N__25813\,
            I => \dataRead7_1\
        );

    \I__5020\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25803\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__25803\,
            I => \N__25792\
        );

    \I__5018\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25789\
        );

    \I__5017\ : InMux
    port map (
            O => \N__25801\,
            I => \N__25786\
        );

    \I__5016\ : InMux
    port map (
            O => \N__25800\,
            I => \N__25779\
        );

    \I__5015\ : InMux
    port map (
            O => \N__25799\,
            I => \N__25779\
        );

    \I__5014\ : InMux
    port map (
            O => \N__25798\,
            I => \N__25779\
        );

    \I__5013\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25773\
        );

    \I__5012\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25773\
        );

    \I__5011\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25769\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__25792\,
            I => \N__25764\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__25789\,
            I => \N__25764\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__25786\,
            I => \N__25761\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__25779\,
            I => \N__25758\
        );

    \I__5006\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25753\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__25773\,
            I => \N__25750\
        );

    \I__5004\ : InMux
    port map (
            O => \N__25772\,
            I => \N__25747\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__25769\,
            I => \N__25744\
        );

    \I__5002\ : Span4Mux_v
    port map (
            O => \N__25764\,
            I => \N__25739\
        );

    \I__5001\ : Span4Mux_h
    port map (
            O => \N__25761\,
            I => \N__25739\
        );

    \I__5000\ : Span4Mux_h
    port map (
            O => \N__25758\,
            I => \N__25736\
        );

    \I__4999\ : CascadeMux
    port map (
            O => \N__25757\,
            I => \N__25717\
        );

    \I__4998\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25712\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__25753\,
            I => \N__25707\
        );

    \I__4996\ : Span4Mux_h
    port map (
            O => \N__25750\,
            I => \N__25707\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__25747\,
            I => \N__25702\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__25744\,
            I => \N__25702\
        );

    \I__4993\ : Span4Mux_h
    port map (
            O => \N__25739\,
            I => \N__25697\
        );

    \I__4992\ : Span4Mux_h
    port map (
            O => \N__25736\,
            I => \N__25697\
        );

    \I__4991\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25680\
        );

    \I__4990\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25680\
        );

    \I__4989\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25680\
        );

    \I__4988\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25680\
        );

    \I__4987\ : InMux
    port map (
            O => \N__25731\,
            I => \N__25680\
        );

    \I__4986\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25680\
        );

    \I__4985\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25680\
        );

    \I__4984\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25680\
        );

    \I__4983\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25669\
        );

    \I__4982\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25669\
        );

    \I__4981\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25669\
        );

    \I__4980\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25669\
        );

    \I__4979\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25669\
        );

    \I__4978\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25656\
        );

    \I__4977\ : InMux
    port map (
            O => \N__25721\,
            I => \N__25656\
        );

    \I__4976\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25656\
        );

    \I__4975\ : InMux
    port map (
            O => \N__25717\,
            I => \N__25656\
        );

    \I__4974\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25656\
        );

    \I__4973\ : InMux
    port map (
            O => \N__25715\,
            I => \N__25656\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__25712\,
            I => \quadWriteZ0Z_5\
        );

    \I__4971\ : Odrv4
    port map (
            O => \N__25707\,
            I => \quadWriteZ0Z_5\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__25702\,
            I => \quadWriteZ0Z_5\
        );

    \I__4969\ : Odrv4
    port map (
            O => \N__25697\,
            I => \quadWriteZ0Z_5\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__25680\,
            I => \quadWriteZ0Z_5\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__25669\,
            I => \quadWriteZ0Z_5\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__25656\,
            I => \quadWriteZ0Z_5\
        );

    \I__4965\ : InMux
    port map (
            O => \N__25641\,
            I => \N__25638\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__25638\,
            I => \N__25635\
        );

    \I__4963\ : Span4Mux_h
    port map (
            O => \N__25635\,
            I => \N__25632\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__25632\,
            I => \N__25629\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__25629\,
            I => \QuadInstance5.Quad_RNO_0_5_3\
        );

    \I__4960\ : IoInMux
    port map (
            O => \N__25626\,
            I => \N__25623\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__25623\,
            I => \N__25620\
        );

    \I__4958\ : Span4Mux_s3_v
    port map (
            O => \N__25620\,
            I => \N__25617\
        );

    \I__4957\ : Span4Mux_v
    port map (
            O => \N__25617\,
            I => \N__25614\
        );

    \I__4956\ : Span4Mux_v
    port map (
            O => \N__25614\,
            I => \N__25611\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__25611\,
            I => \GB_BUFFER_RST_c_i_g_THRU_CO\
        );

    \I__4954\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25604\
        );

    \I__4953\ : InMux
    port map (
            O => \N__25607\,
            I => \N__25601\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__25604\,
            I => \N__25598\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__25601\,
            I => \N__25594\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__25598\,
            I => \N__25591\
        );

    \I__4949\ : CascadeMux
    port map (
            O => \N__25597\,
            I => \N__25588\
        );

    \I__4948\ : Span4Mux_h
    port map (
            O => \N__25594\,
            I => \N__25583\
        );

    \I__4947\ : Span4Mux_v
    port map (
            O => \N__25591\,
            I => \N__25583\
        );

    \I__4946\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25580\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__25583\,
            I => \dataRead5_7\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__25580\,
            I => \dataRead5_7\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__25575\,
            I => \N__25572\
        );

    \I__4942\ : InMux
    port map (
            O => \N__25572\,
            I => \N__25569\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__25569\,
            I => \N__25564\
        );

    \I__4940\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25561\
        );

    \I__4939\ : InMux
    port map (
            O => \N__25567\,
            I => \N__25558\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__25564\,
            I => \N__25555\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__25561\,
            I => \N__25550\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__25558\,
            I => \N__25550\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__25555\,
            I => \dataRead1_7\
        );

    \I__4934\ : Odrv12
    port map (
            O => \N__25550\,
            I => \dataRead1_7\
        );

    \I__4933\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25541\
        );

    \I__4932\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25538\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__25541\,
            I => \N__25535\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__25538\,
            I => \N__25532\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__25535\,
            I => \N__25526\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__25532\,
            I => \N__25526\
        );

    \I__4927\ : InMux
    port map (
            O => \N__25531\,
            I => \N__25523\
        );

    \I__4926\ : Odrv4
    port map (
            O => \N__25526\,
            I => \dataRead1_9\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__25523\,
            I => \dataRead1_9\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__25518\,
            I => \N__25515\
        );

    \I__4923\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25511\
        );

    \I__4922\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25508\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__25511\,
            I => \N__25504\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__25508\,
            I => \N__25501\
        );

    \I__4919\ : InMux
    port map (
            O => \N__25507\,
            I => \N__25498\
        );

    \I__4918\ : Span4Mux_h
    port map (
            O => \N__25504\,
            I => \N__25495\
        );

    \I__4917\ : Span4Mux_v
    port map (
            O => \N__25501\,
            I => \N__25490\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__25498\,
            I => \N__25490\
        );

    \I__4915\ : Odrv4
    port map (
            O => \N__25495\,
            I => \dataRead5_9\
        );

    \I__4914\ : Odrv4
    port map (
            O => \N__25490\,
            I => \dataRead5_9\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__25485\,
            I => \OutReg_ess_RNO_2Z0Z_9_cascade_\
        );

    \I__4912\ : InMux
    port map (
            O => \N__25482\,
            I => \N__25477\
        );

    \I__4911\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25474\
        );

    \I__4910\ : InMux
    port map (
            O => \N__25480\,
            I => \N__25471\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__25477\,
            I => \N__25468\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__25474\,
            I => \N__25463\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__25471\,
            I => \N__25463\
        );

    \I__4906\ : Span4Mux_h
    port map (
            O => \N__25468\,
            I => \N__25460\
        );

    \I__4905\ : Span4Mux_v
    port map (
            O => \N__25463\,
            I => \N__25455\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__25460\,
            I => \N__25455\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__25455\,
            I => \dataRead3_9\
        );

    \I__4902\ : CascadeMux
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__4901\ : InMux
    port map (
            O => \N__25449\,
            I => \N__25446\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__25446\,
            I => \N__25443\
        );

    \I__4899\ : Span4Mux_v
    port map (
            O => \N__25443\,
            I => \N__25439\
        );

    \I__4898\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25435\
        );

    \I__4897\ : Span4Mux_h
    port map (
            O => \N__25439\,
            I => \N__25432\
        );

    \I__4896\ : InMux
    port map (
            O => \N__25438\,
            I => \N__25429\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__25435\,
            I => \N__25424\
        );

    \I__4894\ : Span4Mux_h
    port map (
            O => \N__25432\,
            I => \N__25424\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__25429\,
            I => \dataRead2_9\
        );

    \I__4892\ : Odrv4
    port map (
            O => \N__25424\,
            I => \dataRead2_9\
        );

    \I__4891\ : InMux
    port map (
            O => \N__25419\,
            I => \N__25415\
        );

    \I__4890\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25411\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__25415\,
            I => \N__25408\
        );

    \I__4888\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25405\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__25411\,
            I => \N__25400\
        );

    \I__4886\ : Span4Mux_h
    port map (
            O => \N__25408\,
            I => \N__25400\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__25405\,
            I => \N__25397\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__25400\,
            I => \dataRead6_9\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__25397\,
            I => \dataRead6_9\
        );

    \I__4882\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25388\
        );

    \I__4881\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25384\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__25388\,
            I => \N__25381\
        );

    \I__4879\ : InMux
    port map (
            O => \N__25387\,
            I => \N__25378\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__25384\,
            I => \N__25375\
        );

    \I__4877\ : Span4Mux_h
    port map (
            O => \N__25381\,
            I => \N__25370\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__25378\,
            I => \N__25370\
        );

    \I__4875\ : Span12Mux_v
    port map (
            O => \N__25375\,
            I => \N__25367\
        );

    \I__4874\ : Span4Mux_v
    port map (
            O => \N__25370\,
            I => \N__25364\
        );

    \I__4873\ : Odrv12
    port map (
            O => \N__25367\,
            I => \dataRead7_9\
        );

    \I__4872\ : Odrv4
    port map (
            O => \N__25364\,
            I => \dataRead7_9\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__25359\,
            I => \OutReg_0_4_i_m3_ns_1_9_cascade_\
        );

    \I__4870\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__25353\,
            I => \OutReg_ess_RNO_1Z0Z_9\
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__25350\,
            I => \N__25345\
        );

    \I__4867\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25342\
        );

    \I__4866\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25339\
        );

    \I__4865\ : InMux
    port map (
            O => \N__25345\,
            I => \N__25336\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__25342\,
            I => \N__25331\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__25339\,
            I => \N__25331\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__25336\,
            I => \N__25328\
        );

    \I__4861\ : Span4Mux_v
    port map (
            O => \N__25331\,
            I => \N__25323\
        );

    \I__4860\ : Span4Mux_v
    port map (
            O => \N__25328\,
            I => \N__25323\
        );

    \I__4859\ : Span4Mux_h
    port map (
            O => \N__25323\,
            I => \N__25320\
        );

    \I__4858\ : Odrv4
    port map (
            O => \N__25320\,
            I => \dataRead4_9\
        );

    \I__4857\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25314\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__25314\,
            I => \OutReg_0_5_i_m3_ns_1_9\
        );

    \I__4855\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25307\
        );

    \I__4854\ : InMux
    port map (
            O => \N__25310\,
            I => \N__25304\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__25307\,
            I => \N__25300\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__25304\,
            I => \N__25297\
        );

    \I__4851\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25294\
        );

    \I__4850\ : Span4Mux_v
    port map (
            O => \N__25300\,
            I => \N__25291\
        );

    \I__4849\ : Span4Mux_h
    port map (
            O => \N__25297\,
            I => \N__25286\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__25294\,
            I => \N__25286\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__25291\,
            I => \dataRead1_6\
        );

    \I__4846\ : Odrv4
    port map (
            O => \N__25286\,
            I => \dataRead1_6\
        );

    \I__4845\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25277\
        );

    \I__4844\ : InMux
    port map (
            O => \N__25280\,
            I => \N__25274\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__25277\,
            I => \N__25271\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__25274\,
            I => \N__25268\
        );

    \I__4841\ : Span4Mux_h
    port map (
            O => \N__25271\,
            I => \N__25262\
        );

    \I__4840\ : Span4Mux_h
    port map (
            O => \N__25268\,
            I => \N__25262\
        );

    \I__4839\ : InMux
    port map (
            O => \N__25267\,
            I => \N__25259\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__25262\,
            I => \dataRead5_6\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__25259\,
            I => \dataRead5_6\
        );

    \I__4836\ : CascadeMux
    port map (
            O => \N__25254\,
            I => \OutReg_0_5_i_m3_ns_1_6_cascade_\
        );

    \I__4835\ : CascadeMux
    port map (
            O => \N__25251\,
            I => \N__25248\
        );

    \I__4834\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25245\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__25245\,
            I => \N__25242\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__25242\,
            I => \QuadInstance4.Quad_RNIO30S1Z0Z_9\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__25239\,
            I => \N__25236\
        );

    \I__4830\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25233\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__25233\,
            I => \N__25230\
        );

    \I__4828\ : Span4Mux_s2_v
    port map (
            O => \N__25230\,
            I => \N__25227\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__25227\,
            I => \QuadInstance4.Quad_RNIM10S1Z0Z_7\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__25224\,
            I => \N__25221\
        );

    \I__4825\ : InMux
    port map (
            O => \N__25221\,
            I => \N__25218\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__25218\,
            I => \N__25215\
        );

    \I__4823\ : Span4Mux_h
    port map (
            O => \N__25215\,
            I => \N__25211\
        );

    \I__4822\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25208\
        );

    \I__4821\ : Span4Mux_h
    port map (
            O => \N__25211\,
            I => \N__25205\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__25208\,
            I => \N__25202\
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__25205\,
            I => \dataRead4_15\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__25202\,
            I => \dataRead4_15\
        );

    \I__4817\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25194\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__25194\,
            I => \N__25191\
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__25191\,
            I => \OutReg_0_5_i_m3_ns_1_15\
        );

    \I__4814\ : InMux
    port map (
            O => \N__25188\,
            I => \QuadInstance4.un1_Quad_cry_13\
        );

    \I__4813\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25182\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__4811\ : Span4Mux_v
    port map (
            O => \N__25179\,
            I => \N__25176\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__25176\,
            I => \N__25173\
        );

    \I__4809\ : Odrv4
    port map (
            O => \N__25173\,
            I => \QuadInstance4.un1_Quad_axb_15\
        );

    \I__4808\ : InMux
    port map (
            O => \N__25170\,
            I => \QuadInstance4.un1_Quad_cry_14\
        );

    \I__4807\ : InMux
    port map (
            O => \N__25167\,
            I => \N__25164\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__25164\,
            I => \N__25161\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__25161\,
            I => \QuadInstance4.Quad_RNO_0_4_6\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__25158\,
            I => \N__25155\
        );

    \I__4803\ : InMux
    port map (
            O => \N__25155\,
            I => \N__25152\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__25152\,
            I => \N__25149\
        );

    \I__4801\ : Odrv4
    port map (
            O => \N__25149\,
            I => \QuadInstance4.Quad_RNIL00S1Z0Z_6\
        );

    \I__4800\ : CascadeMux
    port map (
            O => \N__25146\,
            I => \N__25143\
        );

    \I__4799\ : InMux
    port map (
            O => \N__25143\,
            I => \N__25140\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__25140\,
            I => \QuadInstance4.Quad_RNI06TL1Z0Z_10\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__25137\,
            I => \N__25134\
        );

    \I__4796\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25131\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__25131\,
            I => \QuadInstance4.Quad_RNI17TL1Z0Z_11\
        );

    \I__4794\ : InMux
    port map (
            O => \N__25128\,
            I => \N__25125\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__25125\,
            I => \QuadInstance4.Quad_RNO_0_4_11\
        );

    \I__4792\ : CascadeMux
    port map (
            O => \N__25122\,
            I => \N__25119\
        );

    \I__4791\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25116\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__25116\,
            I => \N__25112\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__25115\,
            I => \N__25109\
        );

    \I__4788\ : Span4Mux_v
    port map (
            O => \N__25112\,
            I => \N__25105\
        );

    \I__4787\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25102\
        );

    \I__4786\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25099\
        );

    \I__4785\ : Span4Mux_h
    port map (
            O => \N__25105\,
            I => \N__25096\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__25102\,
            I => \dataRead4_11\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__25099\,
            I => \dataRead4_11\
        );

    \I__4782\ : Odrv4
    port map (
            O => \N__25096\,
            I => \dataRead4_11\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__25089\,
            I => \N__25084\
        );

    \I__4780\ : CascadeMux
    port map (
            O => \N__25088\,
            I => \N__25081\
        );

    \I__4779\ : InMux
    port map (
            O => \N__25087\,
            I => \N__25078\
        );

    \I__4778\ : InMux
    port map (
            O => \N__25084\,
            I => \N__25075\
        );

    \I__4777\ : InMux
    port map (
            O => \N__25081\,
            I => \N__25072\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__25078\,
            I => \N__25069\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__25075\,
            I => \dataRead4_6\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__25072\,
            I => \dataRead4_6\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__25069\,
            I => \dataRead4_6\
        );

    \I__4772\ : InMux
    port map (
            O => \N__25062\,
            I => \QuadInstance4.un1_Quad_cry_4\
        );

    \I__4771\ : InMux
    port map (
            O => \N__25059\,
            I => \QuadInstance4.un1_Quad_cry_5\
        );

    \I__4770\ : InMux
    port map (
            O => \N__25056\,
            I => \QuadInstance4.un1_Quad_cry_6\
        );

    \I__4769\ : InMux
    port map (
            O => \N__25053\,
            I => \bfn_15_4_0_\
        );

    \I__4768\ : InMux
    port map (
            O => \N__25050\,
            I => \N__25047\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__25047\,
            I => \N__25044\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__25044\,
            I => \N__25041\
        );

    \I__4765\ : Span4Mux_h
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__25038\,
            I => \QuadInstance4.Quad_RNO_0_4_9\
        );

    \I__4763\ : InMux
    port map (
            O => \N__25035\,
            I => \QuadInstance4.un1_Quad_cry_8\
        );

    \I__4762\ : InMux
    port map (
            O => \N__25032\,
            I => \QuadInstance4.un1_Quad_cry_9\
        );

    \I__4761\ : InMux
    port map (
            O => \N__25029\,
            I => \QuadInstance4.un1_Quad_cry_10\
        );

    \I__4760\ : InMux
    port map (
            O => \N__25026\,
            I => \QuadInstance4.un1_Quad_cry_11\
        );

    \I__4759\ : InMux
    port map (
            O => \N__25023\,
            I => \QuadInstance4.un1_Quad_cry_12\
        );

    \I__4758\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25017\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__25017\,
            I => \N__25014\
        );

    \I__4756\ : Span4Mux_s3_v
    port map (
            O => \N__25014\,
            I => \N__25011\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__25011\,
            I => \N__25008\
        );

    \I__4754\ : Span4Mux_v
    port map (
            O => \N__25008\,
            I => \N__25005\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__25005\,
            I => \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_3\
        );

    \I__4752\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24999\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__24999\,
            I => \N__24996\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__24996\,
            I => \N__24993\
        );

    \I__4749\ : Sp12to4
    port map (
            O => \N__24993\,
            I => \N__24990\
        );

    \I__4748\ : Span12Mux_s6_v
    port map (
            O => \N__24990\,
            I => \N__24987\
        );

    \I__4747\ : Odrv12
    port map (
            O => \N__24987\,
            I => \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_3\
        );

    \I__4746\ : InMux
    port map (
            O => \N__24984\,
            I => \bfn_15_2_0_\
        );

    \I__4745\ : IoInMux
    port map (
            O => \N__24981\,
            I => \N__24978\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__24978\,
            I => \N__24975\
        );

    \I__4743\ : IoSpan4Mux
    port map (
            O => \N__24975\,
            I => \N__24972\
        );

    \I__4742\ : Span4Mux_s2_v
    port map (
            O => \N__24972\,
            I => \N__24969\
        );

    \I__4741\ : Span4Mux_v
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__4740\ : Sp12to4
    port map (
            O => \N__24966\,
            I => \N__24963\
        );

    \I__4739\ : Span12Mux_v
    port map (
            O => \N__24963\,
            I => \N__24959\
        );

    \I__4738\ : InMux
    port map (
            O => \N__24962\,
            I => \N__24956\
        );

    \I__4737\ : Odrv12
    port map (
            O => \N__24959\,
            I => \PWM4_c\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__24956\,
            I => \PWM4_c\
        );

    \I__4735\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24948\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__24948\,
            I => \N__24945\
        );

    \I__4733\ : Span4Mux_h
    port map (
            O => \N__24945\,
            I => \N__24942\
        );

    \I__4732\ : Odrv4
    port map (
            O => \N__24942\,
            I => \QuadInstance4.Quad_RNO_0_3_1\
        );

    \I__4731\ : InMux
    port map (
            O => \N__24939\,
            I => \QuadInstance4.un1_Quad_cry_0\
        );

    \I__4730\ : InMux
    port map (
            O => \N__24936\,
            I => \QuadInstance4.un1_Quad_cry_1\
        );

    \I__4729\ : InMux
    port map (
            O => \N__24933\,
            I => \QuadInstance4.un1_Quad_cry_2\
        );

    \I__4728\ : InMux
    port map (
            O => \N__24930\,
            I => \N__24927\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__24927\,
            I => \N__24924\
        );

    \I__4726\ : Span4Mux_h
    port map (
            O => \N__24924\,
            I => \N__24921\
        );

    \I__4725\ : Odrv4
    port map (
            O => \N__24921\,
            I => \QuadInstance4.Quad_RNO_0_4_4\
        );

    \I__4724\ : InMux
    port map (
            O => \N__24918\,
            I => \QuadInstance4.un1_Quad_cry_3\
        );

    \I__4723\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24911\
        );

    \I__4722\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24907\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__24911\,
            I => \N__24904\
        );

    \I__4720\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24901\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__24907\,
            I => \PWMInstance4.periodCounterZ0Z_14\
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__24904\,
            I => \PWMInstance4.periodCounterZ0Z_14\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__24901\,
            I => \PWMInstance4.periodCounterZ0Z_14\
        );

    \I__4716\ : InMux
    port map (
            O => \N__24894\,
            I => \PWMInstance4.un1_periodCounter_2_cry_13\
        );

    \I__4715\ : InMux
    port map (
            O => \N__24891\,
            I => \PWMInstance4.un1_periodCounter_2_cry_14\
        );

    \I__4714\ : InMux
    port map (
            O => \N__24888\,
            I => \bfn_14_18_0_\
        );

    \I__4713\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24882\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__24882\,
            I => \N__24879\
        );

    \I__4711\ : Span4Mux_s2_v
    port map (
            O => \N__24879\,
            I => \N__24876\
        );

    \I__4710\ : Span4Mux_v
    port map (
            O => \N__24876\,
            I => \N__24873\
        );

    \I__4709\ : Span4Mux_v
    port map (
            O => \N__24873\,
            I => \N__24870\
        );

    \I__4708\ : Odrv4
    port map (
            O => \N__24870\,
            I => \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_3\
        );

    \I__4707\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24864\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__4705\ : Span12Mux_h
    port map (
            O => \N__24861\,
            I => \N__24858\
        );

    \I__4704\ : Span12Mux_v
    port map (
            O => \N__24858\,
            I => \N__24855\
        );

    \I__4703\ : Odrv12
    port map (
            O => \N__24855\,
            I => \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_3\
        );

    \I__4702\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24849\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24846\
        );

    \I__4700\ : Span4Mux_h
    port map (
            O => \N__24846\,
            I => \N__24843\
        );

    \I__4699\ : Sp12to4
    port map (
            O => \N__24843\,
            I => \N__24840\
        );

    \I__4698\ : Span12Mux_s9_v
    port map (
            O => \N__24840\,
            I => \N__24837\
        );

    \I__4697\ : Odrv12
    port map (
            O => \N__24837\,
            I => \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_3\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__24834\,
            I => \N__24829\
        );

    \I__4695\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24826\
        );

    \I__4694\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24823\
        );

    \I__4693\ : InMux
    port map (
            O => \N__24829\,
            I => \N__24820\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__24826\,
            I => \PWMInstance4.periodCounterZ0Z_5\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__24823\,
            I => \PWMInstance4.periodCounterZ0Z_5\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__24820\,
            I => \PWMInstance4.periodCounterZ0Z_5\
        );

    \I__4689\ : InMux
    port map (
            O => \N__24813\,
            I => \PWMInstance4.un1_periodCounter_2_cry_4\
        );

    \I__4688\ : InMux
    port map (
            O => \N__24810\,
            I => \PWMInstance4.un1_periodCounter_2_cry_5\
        );

    \I__4687\ : InMux
    port map (
            O => \N__24807\,
            I => \PWMInstance4.un1_periodCounter_2_cry_6\
        );

    \I__4686\ : InMux
    port map (
            O => \N__24804\,
            I => \bfn_14_17_0_\
        );

    \I__4685\ : InMux
    port map (
            O => \N__24801\,
            I => \PWMInstance4.un1_periodCounter_2_cry_8\
        );

    \I__4684\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24793\
        );

    \I__4683\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24788\
        );

    \I__4682\ : InMux
    port map (
            O => \N__24796\,
            I => \N__24788\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__24793\,
            I => \PWMInstance4.periodCounterZ0Z_10\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__24788\,
            I => \PWMInstance4.periodCounterZ0Z_10\
        );

    \I__4679\ : InMux
    port map (
            O => \N__24783\,
            I => \PWMInstance4.un1_periodCounter_2_cry_9\
        );

    \I__4678\ : CascadeMux
    port map (
            O => \N__24780\,
            I => \N__24777\
        );

    \I__4677\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24772\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__24776\,
            I => \N__24769\
        );

    \I__4675\ : InMux
    port map (
            O => \N__24775\,
            I => \N__24766\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__24772\,
            I => \N__24763\
        );

    \I__4673\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24760\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__24766\,
            I => \PWMInstance4.periodCounterZ0Z_11\
        );

    \I__4671\ : Odrv4
    port map (
            O => \N__24763\,
            I => \PWMInstance4.periodCounterZ0Z_11\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__24760\,
            I => \PWMInstance4.periodCounterZ0Z_11\
        );

    \I__4669\ : InMux
    port map (
            O => \N__24753\,
            I => \PWMInstance4.un1_periodCounter_2_cry_10\
        );

    \I__4668\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24746\
        );

    \I__4667\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24742\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__24746\,
            I => \N__24739\
        );

    \I__4665\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24736\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__24742\,
            I => \PWMInstance4.periodCounterZ0Z_12\
        );

    \I__4663\ : Odrv4
    port map (
            O => \N__24739\,
            I => \PWMInstance4.periodCounterZ0Z_12\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__24736\,
            I => \PWMInstance4.periodCounterZ0Z_12\
        );

    \I__4661\ : InMux
    port map (
            O => \N__24729\,
            I => \PWMInstance4.un1_periodCounter_2_cry_11\
        );

    \I__4660\ : InMux
    port map (
            O => \N__24726\,
            I => \PWMInstance4.un1_periodCounter_2_cry_12\
        );

    \I__4659\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24720\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__24720\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_14\
        );

    \I__4657\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24714\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__24714\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_15\
        );

    \I__4655\ : InMux
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__24708\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_12\
        );

    \I__4653\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24702\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__24702\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_13\
        );

    \I__4651\ : InMux
    port map (
            O => \N__24699\,
            I => \PWMInstance4.un1_periodCounter_2_cry_0\
        );

    \I__4650\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24691\
        );

    \I__4649\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24688\
        );

    \I__4648\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24685\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__24691\,
            I => \PWMInstance4.periodCounterZ0Z_2\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__24688\,
            I => \PWMInstance4.periodCounterZ0Z_2\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__24685\,
            I => \PWMInstance4.periodCounterZ0Z_2\
        );

    \I__4644\ : InMux
    port map (
            O => \N__24678\,
            I => \PWMInstance4.un1_periodCounter_2_cry_1\
        );

    \I__4643\ : CascadeMux
    port map (
            O => \N__24675\,
            I => \N__24670\
        );

    \I__4642\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24667\
        );

    \I__4641\ : InMux
    port map (
            O => \N__24673\,
            I => \N__24662\
        );

    \I__4640\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24662\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__24667\,
            I => \PWMInstance4.periodCounterZ0Z_3\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__24662\,
            I => \PWMInstance4.periodCounterZ0Z_3\
        );

    \I__4637\ : InMux
    port map (
            O => \N__24657\,
            I => \PWMInstance4.un1_periodCounter_2_cry_2\
        );

    \I__4636\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24649\
        );

    \I__4635\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24644\
        );

    \I__4634\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24644\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__24649\,
            I => \PWMInstance4.periodCounterZ0Z_4\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__24644\,
            I => \PWMInstance4.periodCounterZ0Z_4\
        );

    \I__4631\ : InMux
    port map (
            O => \N__24639\,
            I => \PWMInstance4.un1_periodCounter_2_cry_3\
        );

    \I__4630\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24629\
        );

    \I__4629\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24629\
        );

    \I__4628\ : InMux
    port map (
            O => \N__24634\,
            I => \N__24626\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__24629\,
            I => \pwmWriteZ0Z_3\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__24626\,
            I => \pwmWriteZ0Z_3\
        );

    \I__4625\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24615\
        );

    \I__4624\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24615\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__24615\,
            I => \pwmWrite_fastZ0Z_3\
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__24612\,
            I => \N__24608\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__24611\,
            I => \N__24605\
        );

    \I__4620\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24594\
        );

    \I__4619\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24594\
        );

    \I__4618\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24594\
        );

    \I__4617\ : InMux
    port map (
            O => \N__24603\,
            I => \N__24594\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__24594\,
            I => \PWMInstance3.clkCountZ0Z_1\
        );

    \I__4615\ : InMux
    port map (
            O => \N__24591\,
            I => \N__24579\
        );

    \I__4614\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24579\
        );

    \I__4613\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24579\
        );

    \I__4612\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24579\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__24579\,
            I => \PWMInstance3.clkCountZ0Z_0\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__24576\,
            I => \PWMInstance3.un1_periodCounter12_1_0_a2_0_6_cascade_\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__24573\,
            I => \PWMInstance3.un1_periodCounter12_1_0_a2_0_14_cascade_\
        );

    \I__4608\ : InMux
    port map (
            O => \N__24570\,
            I => \N__24567\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__24567\,
            I => \N__24564\
        );

    \I__4606\ : Span4Mux_v
    port map (
            O => \N__24564\,
            I => \N__24561\
        );

    \I__4605\ : Odrv4
    port map (
            O => \N__24561\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_9\
        );

    \I__4604\ : CEMux
    port map (
            O => \N__24558\,
            I => \N__24553\
        );

    \I__4603\ : CEMux
    port map (
            O => \N__24557\,
            I => \N__24549\
        );

    \I__4602\ : CEMux
    port map (
            O => \N__24556\,
            I => \N__24546\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__24553\,
            I => \N__24543\
        );

    \I__4600\ : CEMux
    port map (
            O => \N__24552\,
            I => \N__24540\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__24549\,
            I => \N__24536\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__24546\,
            I => \N__24533\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__24543\,
            I => \N__24530\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__24540\,
            I => \N__24527\
        );

    \I__4595\ : CEMux
    port map (
            O => \N__24539\,
            I => \N__24524\
        );

    \I__4594\ : Span4Mux_v
    port map (
            O => \N__24536\,
            I => \N__24521\
        );

    \I__4593\ : Span4Mux_h
    port map (
            O => \N__24533\,
            I => \N__24518\
        );

    \I__4592\ : Span4Mux_h
    port map (
            O => \N__24530\,
            I => \N__24513\
        );

    \I__4591\ : Span4Mux_h
    port map (
            O => \N__24527\,
            I => \N__24513\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__24524\,
            I => \N__24510\
        );

    \I__4589\ : Span4Mux_h
    port map (
            O => \N__24521\,
            I => \N__24507\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__24518\,
            I => \PWMInstance6.pwmWrite_0_6\
        );

    \I__4587\ : Odrv4
    port map (
            O => \N__24513\,
            I => \PWMInstance6.pwmWrite_0_6\
        );

    \I__4586\ : Odrv12
    port map (
            O => \N__24510\,
            I => \PWMInstance6.pwmWrite_0_6\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__24507\,
            I => \PWMInstance6.pwmWrite_0_6\
        );

    \I__4584\ : InMux
    port map (
            O => \N__24498\,
            I => \N__24495\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__24495\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_3\
        );

    \I__4582\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24489\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__24489\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_2\
        );

    \I__4580\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24482\
        );

    \I__4579\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24479\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__24482\,
            I => \data_receivedZ0Z_8\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__24479\,
            I => \data_receivedZ0Z_8\
        );

    \I__4576\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24470\
        );

    \I__4575\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24467\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__24470\,
            I => \data_receivedZ0Z_9\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__24467\,
            I => \data_receivedZ0Z_9\
        );

    \I__4572\ : CEMux
    port map (
            O => \N__24462\,
            I => \N__24458\
        );

    \I__4571\ : CEMux
    port map (
            O => \N__24461\,
            I => \N__24455\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__24458\,
            I => \N_870_i\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__24455\,
            I => \N_870_i\
        );

    \I__4568\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24446\
        );

    \I__4567\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24443\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__24446\,
            I => \data_receivedZ0Z_5\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__24443\,
            I => \data_receivedZ0Z_5\
        );

    \I__4564\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24434\
        );

    \I__4563\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24431\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__24434\,
            I => \data_receivedZ0Z_6\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__24431\,
            I => \data_receivedZ0Z_6\
        );

    \I__4560\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24422\
        );

    \I__4559\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24419\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__24422\,
            I => \data_receivedZ0Z_7\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__24419\,
            I => \data_receivedZ0Z_7\
        );

    \I__4556\ : InMux
    port map (
            O => \N__24414\,
            I => \N__24411\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__24411\,
            I => \N__24407\
        );

    \I__4554\ : InMux
    port map (
            O => \N__24410\,
            I => \N__24403\
        );

    \I__4553\ : Span4Mux_v
    port map (
            O => \N__24407\,
            I => \N__24400\
        );

    \I__4552\ : InMux
    port map (
            O => \N__24406\,
            I => \N__24397\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__24403\,
            I => \N__24394\
        );

    \I__4550\ : Span4Mux_v
    port map (
            O => \N__24400\,
            I => \N__24389\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__24397\,
            I => \N__24389\
        );

    \I__4548\ : Span4Mux_h
    port map (
            O => \N__24394\,
            I => \N__24386\
        );

    \I__4547\ : Span4Mux_h
    port map (
            O => \N__24389\,
            I => \N__24383\
        );

    \I__4546\ : Span4Mux_v
    port map (
            O => \N__24386\,
            I => \N__24380\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__24383\,
            I => \dataRead2_3\
        );

    \I__4544\ : Odrv4
    port map (
            O => \N__24380\,
            I => \dataRead2_3\
        );

    \I__4543\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24371\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__24374\,
            I => \N__24368\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__24371\,
            I => \N__24364\
        );

    \I__4540\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24361\
        );

    \I__4539\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24358\
        );

    \I__4538\ : Span4Mux_h
    port map (
            O => \N__24364\,
            I => \N__24355\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__24361\,
            I => \N__24352\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__24358\,
            I => \N__24349\
        );

    \I__4535\ : Span4Mux_v
    port map (
            O => \N__24355\,
            I => \N__24346\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__24352\,
            I => \N__24341\
        );

    \I__4533\ : Span4Mux_h
    port map (
            O => \N__24349\,
            I => \N__24341\
        );

    \I__4532\ : Odrv4
    port map (
            O => \N__24346\,
            I => \dataRead3_3\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__24341\,
            I => \dataRead3_3\
        );

    \I__4530\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24332\
        );

    \I__4529\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24329\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__24332\,
            I => \N__24326\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24323\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__24326\,
            I => \N__24320\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__24323\,
            I => \dataRead3_15\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__24320\,
            I => \dataRead3_15\
        );

    \I__4523\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24311\
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__24314\,
            I => \N__24308\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__24311\,
            I => \N__24305\
        );

    \I__4520\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24302\
        );

    \I__4519\ : Span4Mux_h
    port map (
            O => \N__24305\,
            I => \N__24299\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24294\
        );

    \I__4517\ : Span4Mux_h
    port map (
            O => \N__24299\,
            I => \N__24294\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__24294\,
            I => \dataRead2_15\
        );

    \I__4515\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24287\
        );

    \I__4514\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24284\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__24287\,
            I => \N__24281\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__24284\,
            I => \N__24276\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__24281\,
            I => \N__24276\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__24276\,
            I => \dataRead7_15\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__24273\,
            I => \N__24270\
        );

    \I__4508\ : InMux
    port map (
            O => \N__24270\,
            I => \N__24266\
        );

    \I__4507\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24263\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__24266\,
            I => \N__24260\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__24263\,
            I => \N__24257\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__24260\,
            I => \N__24252\
        );

    \I__4503\ : Span4Mux_h
    port map (
            O => \N__24257\,
            I => \N__24252\
        );

    \I__4502\ : Odrv4
    port map (
            O => \N__24252\,
            I => \dataRead6_15\
        );

    \I__4501\ : CascadeMux
    port map (
            O => \N__24249\,
            I => \OutReg_0_4_i_m3_ns_1_15_cascade_\
        );

    \I__4500\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24243\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__24243\,
            I => \N__24239\
        );

    \I__4498\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24236\
        );

    \I__4497\ : Span4Mux_h
    port map (
            O => \N__24239\,
            I => \N__24233\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__24236\,
            I => \dataRead5_15\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__24233\,
            I => \dataRead5_15\
        );

    \I__4494\ : CascadeMux
    port map (
            O => \N__24228\,
            I => \N__24224\
        );

    \I__4493\ : InMux
    port map (
            O => \N__24227\,
            I => \N__24221\
        );

    \I__4492\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24218\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__24221\,
            I => \N__24213\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__24218\,
            I => \N__24213\
        );

    \I__4489\ : Odrv4
    port map (
            O => \N__24213\,
            I => \dataRead1_15\
        );

    \I__4488\ : CascadeMux
    port map (
            O => \N__24210\,
            I => \N__24205\
        );

    \I__4487\ : CascadeMux
    port map (
            O => \N__24209\,
            I => \N__24202\
        );

    \I__4486\ : InMux
    port map (
            O => \N__24208\,
            I => \N__24183\
        );

    \I__4485\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24183\
        );

    \I__4484\ : InMux
    port map (
            O => \N__24202\,
            I => \N__24183\
        );

    \I__4483\ : InMux
    port map (
            O => \N__24201\,
            I => \N__24183\
        );

    \I__4482\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24183\
        );

    \I__4481\ : InMux
    port map (
            O => \N__24199\,
            I => \N__24183\
        );

    \I__4480\ : CascadeMux
    port map (
            O => \N__24198\,
            I => \N__24175\
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__24197\,
            I => \N__24170\
        );

    \I__4478\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24167\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__24183\,
            I => \N__24164\
        );

    \I__4476\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24157\
        );

    \I__4475\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24157\
        );

    \I__4474\ : InMux
    port map (
            O => \N__24180\,
            I => \N__24157\
        );

    \I__4473\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24144\
        );

    \I__4472\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24144\
        );

    \I__4471\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24144\
        );

    \I__4470\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24144\
        );

    \I__4469\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24144\
        );

    \I__4468\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24144\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__24167\,
            I => \QuadInstance1.count_enable\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__24164\,
            I => \QuadInstance1.count_enable\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__24157\,
            I => \QuadInstance1.count_enable\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__24144\,
            I => \QuadInstance1.count_enable\
        );

    \I__4463\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24132\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__24132\,
            I => \QuadInstance1.Quad_RNO_0_1_12\
        );

    \I__4461\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24125\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__24128\,
            I => \N__24122\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__24125\,
            I => \N__24118\
        );

    \I__4458\ : InMux
    port map (
            O => \N__24122\,
            I => \N__24115\
        );

    \I__4457\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24112\
        );

    \I__4456\ : Span4Mux_v
    port map (
            O => \N__24118\,
            I => \N__24109\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__24115\,
            I => \dataRead1_12\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__24112\,
            I => \dataRead1_12\
        );

    \I__4453\ : Odrv4
    port map (
            O => \N__24109\,
            I => \dataRead1_12\
        );

    \I__4452\ : InMux
    port map (
            O => \N__24102\,
            I => \N__24092\
        );

    \I__4451\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24087\
        );

    \I__4450\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24087\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__24099\,
            I => \N__24081\
        );

    \I__4448\ : InMux
    port map (
            O => \N__24098\,
            I => \N__24077\
        );

    \I__4447\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24072\
        );

    \I__4446\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24072\
        );

    \I__4445\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24069\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__24092\,
            I => \N__24066\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__24087\,
            I => \N__24063\
        );

    \I__4442\ : InMux
    port map (
            O => \N__24086\,
            I => \N__24060\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__24085\,
            I => \N__24056\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__24084\,
            I => \N__24053\
        );

    \I__4439\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24045\
        );

    \I__4438\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24045\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__24077\,
            I => \N__24042\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__24072\,
            I => \N__24037\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__24069\,
            I => \N__24037\
        );

    \I__4434\ : Span4Mux_v
    port map (
            O => \N__24066\,
            I => \N__24032\
        );

    \I__4433\ : Span4Mux_v
    port map (
            O => \N__24063\,
            I => \N__24032\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__24060\,
            I => \N__24029\
        );

    \I__4431\ : InMux
    port map (
            O => \N__24059\,
            I => \N__24018\
        );

    \I__4430\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24011\
        );

    \I__4429\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24011\
        );

    \I__4428\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24011\
        );

    \I__4427\ : InMux
    port map (
            O => \N__24051\,
            I => \N__24001\
        );

    \I__4426\ : InMux
    port map (
            O => \N__24050\,
            I => \N__23998\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__24045\,
            I => \N__23993\
        );

    \I__4424\ : Span4Mux_v
    port map (
            O => \N__24042\,
            I => \N__23993\
        );

    \I__4423\ : Span4Mux_h
    port map (
            O => \N__24037\,
            I => \N__23990\
        );

    \I__4422\ : Sp12to4
    port map (
            O => \N__24032\,
            I => \N__23985\
        );

    \I__4421\ : Span12Mux_v
    port map (
            O => \N__24029\,
            I => \N__23985\
        );

    \I__4420\ : InMux
    port map (
            O => \N__24028\,
            I => \N__23968\
        );

    \I__4419\ : InMux
    port map (
            O => \N__24027\,
            I => \N__23968\
        );

    \I__4418\ : InMux
    port map (
            O => \N__24026\,
            I => \N__23968\
        );

    \I__4417\ : InMux
    port map (
            O => \N__24025\,
            I => \N__23968\
        );

    \I__4416\ : InMux
    port map (
            O => \N__24024\,
            I => \N__23968\
        );

    \I__4415\ : InMux
    port map (
            O => \N__24023\,
            I => \N__23968\
        );

    \I__4414\ : InMux
    port map (
            O => \N__24022\,
            I => \N__23968\
        );

    \I__4413\ : InMux
    port map (
            O => \N__24021\,
            I => \N__23968\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__24018\,
            I => \N__23963\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__23963\
        );

    \I__4410\ : InMux
    port map (
            O => \N__24010\,
            I => \N__23950\
        );

    \I__4409\ : InMux
    port map (
            O => \N__24009\,
            I => \N__23950\
        );

    \I__4408\ : InMux
    port map (
            O => \N__24008\,
            I => \N__23950\
        );

    \I__4407\ : InMux
    port map (
            O => \N__24007\,
            I => \N__23950\
        );

    \I__4406\ : InMux
    port map (
            O => \N__24006\,
            I => \N__23950\
        );

    \I__4405\ : InMux
    port map (
            O => \N__24005\,
            I => \N__23950\
        );

    \I__4404\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23947\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__24001\,
            I => \quadWriteZ0Z_1\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__23998\,
            I => \quadWriteZ0Z_1\
        );

    \I__4401\ : Odrv4
    port map (
            O => \N__23993\,
            I => \quadWriteZ0Z_1\
        );

    \I__4400\ : Odrv4
    port map (
            O => \N__23990\,
            I => \quadWriteZ0Z_1\
        );

    \I__4399\ : Odrv12
    port map (
            O => \N__23985\,
            I => \quadWriteZ0Z_1\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__23968\,
            I => \quadWriteZ0Z_1\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__23963\,
            I => \quadWriteZ0Z_1\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__23950\,
            I => \quadWriteZ0Z_1\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__23947\,
            I => \quadWriteZ0Z_1\
        );

    \I__4394\ : InMux
    port map (
            O => \N__23928\,
            I => \N__23925\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__23925\,
            I => \QuadInstance1.Quad_RNO_0_1_13\
        );

    \I__4392\ : InMux
    port map (
            O => \N__23922\,
            I => \N__23919\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__23919\,
            I => \N__23914\
        );

    \I__4390\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23911\
        );

    \I__4389\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23908\
        );

    \I__4388\ : Span4Mux_v
    port map (
            O => \N__23914\,
            I => \N__23905\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__23911\,
            I => \dataRead1_13\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__23908\,
            I => \dataRead1_13\
        );

    \I__4385\ : Odrv4
    port map (
            O => \N__23905\,
            I => \dataRead1_13\
        );

    \I__4384\ : InMux
    port map (
            O => \N__23898\,
            I => \N__23894\
        );

    \I__4383\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23891\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__23894\,
            I => \N__23887\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__23891\,
            I => \N__23884\
        );

    \I__4380\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23881\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__23887\,
            I => \N__23878\
        );

    \I__4378\ : Span4Mux_v
    port map (
            O => \N__23884\,
            I => \N__23873\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__23881\,
            I => \N__23873\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__23878\,
            I => \dataRead1_1\
        );

    \I__4375\ : Odrv4
    port map (
            O => \N__23873\,
            I => \dataRead1_1\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__23868\,
            I => \N__23865\
        );

    \I__4373\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23862\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__23862\,
            I => \N__23859\
        );

    \I__4371\ : Span4Mux_h
    port map (
            O => \N__23859\,
            I => \N__23855\
        );

    \I__4370\ : InMux
    port map (
            O => \N__23858\,
            I => \N__23851\
        );

    \I__4369\ : Span4Mux_h
    port map (
            O => \N__23855\,
            I => \N__23848\
        );

    \I__4368\ : InMux
    port map (
            O => \N__23854\,
            I => \N__23845\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__23851\,
            I => \dataRead5_1\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__23848\,
            I => \dataRead5_1\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__23845\,
            I => \dataRead5_1\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__23838\,
            I => \OutReg_ess_RNO_2Z0Z_1_cascade_\
        );

    \I__4363\ : InMux
    port map (
            O => \N__23835\,
            I => \N__23831\
        );

    \I__4362\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23828\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__23831\,
            I => \N__23822\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__23828\,
            I => \N__23822\
        );

    \I__4359\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23819\
        );

    \I__4358\ : Span12Mux_s7_v
    port map (
            O => \N__23822\,
            I => \N__23816\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__23819\,
            I => \dataRead2_1\
        );

    \I__4356\ : Odrv12
    port map (
            O => \N__23816\,
            I => \dataRead2_1\
        );

    \I__4355\ : InMux
    port map (
            O => \N__23811\,
            I => \N__23808\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__23808\,
            I => \N__23804\
        );

    \I__4353\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23801\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__23804\,
            I => \N__23795\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__23801\,
            I => \N__23795\
        );

    \I__4350\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23792\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__23795\,
            I => \dataRead3_1\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__23792\,
            I => \dataRead3_1\
        );

    \I__4347\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23784\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23779\
        );

    \I__4345\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23776\
        );

    \I__4344\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23773\
        );

    \I__4343\ : Span4Mux_h
    port map (
            O => \N__23779\,
            I => \N__23770\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__23776\,
            I => \N__23767\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__23773\,
            I => \dataRead6_1\
        );

    \I__4340\ : Odrv4
    port map (
            O => \N__23770\,
            I => \dataRead6_1\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__23767\,
            I => \dataRead6_1\
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__23760\,
            I => \OutReg_0_4_i_m3_ns_1_1_cascade_\
        );

    \I__4337\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23754\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__23754\,
            I => \OutReg_ess_RNO_1Z0Z_1\
        );

    \I__4335\ : InMux
    port map (
            O => \N__23751\,
            I => \N__23748\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__23748\,
            I => \OutReg_0_5_i_m3_ns_1_1\
        );

    \I__4333\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23742\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__23742\,
            I => \N__23738\
        );

    \I__4331\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23735\
        );

    \I__4330\ : Span4Mux_h
    port map (
            O => \N__23738\,
            I => \N__23729\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__23735\,
            I => \N__23729\
        );

    \I__4328\ : InMux
    port map (
            O => \N__23734\,
            I => \N__23726\
        );

    \I__4327\ : Span4Mux_v
    port map (
            O => \N__23729\,
            I => \N__23721\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__23726\,
            I => \N__23721\
        );

    \I__4325\ : Odrv4
    port map (
            O => \N__23721\,
            I => \dataRead3_5\
        );

    \I__4324\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23714\
        );

    \I__4323\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23711\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__23714\,
            I => \N__23707\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__23711\,
            I => \N__23704\
        );

    \I__4320\ : InMux
    port map (
            O => \N__23710\,
            I => \N__23701\
        );

    \I__4319\ : Span4Mux_v
    port map (
            O => \N__23707\,
            I => \N__23696\
        );

    \I__4318\ : Span4Mux_h
    port map (
            O => \N__23704\,
            I => \N__23696\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__23701\,
            I => \N__23693\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__23696\,
            I => \N__23688\
        );

    \I__4315\ : Span4Mux_h
    port map (
            O => \N__23693\,
            I => \N__23688\
        );

    \I__4314\ : Odrv4
    port map (
            O => \N__23688\,
            I => \dataRead2_5\
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__4312\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__23679\,
            I => \QuadInstance1.Quad_RNIUN0OZ0Z_7\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__4309\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__23670\,
            I => \QuadInstance1.Quad_RNIPI0OZ0Z_2\
        );

    \I__4307\ : CascadeMux
    port map (
            O => \N__23667\,
            I => \N__23664\
        );

    \I__4306\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23661\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__23661\,
            I => \QuadInstance1.Quad_RNIQJ0OZ0Z_3\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__23658\,
            I => \N__23655\
        );

    \I__4303\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23652\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__23652\,
            I => \QuadInstance1.Quad_RNIAR5DZ0Z_12\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__23649\,
            I => \N__23646\
        );

    \I__4300\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23643\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__23643\,
            I => \QuadInstance1.Quad_RNIBS5DZ0Z_13\
        );

    \I__4298\ : InMux
    port map (
            O => \N__23640\,
            I => \N__23637\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__23637\,
            I => \QuadInstance1.Quad_RNICT5DZ0Z_14\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__23634\,
            I => \N__23631\
        );

    \I__4295\ : InMux
    port map (
            O => \N__23631\,
            I => \N__23628\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__23628\,
            I => \QuadInstance1.Quad_RNIVO0OZ0Z_8\
        );

    \I__4293\ : CascadeMux
    port map (
            O => \N__23625\,
            I => \N__23619\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__23624\,
            I => \N__23615\
        );

    \I__4291\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23599\
        );

    \I__4290\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23599\
        );

    \I__4289\ : InMux
    port map (
            O => \N__23619\,
            I => \N__23599\
        );

    \I__4288\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23599\
        );

    \I__4287\ : InMux
    port map (
            O => \N__23615\,
            I => \N__23599\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__23614\,
            I => \N__23596\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__23613\,
            I => \N__23592\
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__23612\,
            I => \N__23589\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__23611\,
            I => \N__23585\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__23610\,
            I => \N__23582\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__23599\,
            I => \N__23576\
        );

    \I__4280\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23563\
        );

    \I__4279\ : InMux
    port map (
            O => \N__23595\,
            I => \N__23563\
        );

    \I__4278\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23563\
        );

    \I__4277\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23563\
        );

    \I__4276\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23563\
        );

    \I__4275\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23563\
        );

    \I__4274\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23554\
        );

    \I__4273\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23554\
        );

    \I__4272\ : InMux
    port map (
            O => \N__23580\,
            I => \N__23554\
        );

    \I__4271\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23554\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__23576\,
            I => \QuadInstance1.un1_count_enable_i_a2_0_1\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__23563\,
            I => \QuadInstance1.un1_count_enable_i_a2_0_1\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__23554\,
            I => \QuadInstance1.un1_count_enable_i_a2_0_1\
        );

    \I__4267\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23544\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__23544\,
            I => \QuadInstance1.un1_Quad_axb_15\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__23541\,
            I => \QuadInstance1.count_enable_cascade_\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__23538\,
            I => \N__23535\
        );

    \I__4263\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23532\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__23532\,
            I => \QuadInstance1.Quad_RNIOH0OZ0Z_1\
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__23529\,
            I => \N__23526\
        );

    \I__4260\ : InMux
    port map (
            O => \N__23526\,
            I => \N__23523\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__23523\,
            I => \QuadInstance1.Quad_RNITM0OZ0Z_6\
        );

    \I__4258\ : CascadeMux
    port map (
            O => \N__23520\,
            I => \N__23517\
        );

    \I__4257\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23514\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__23514\,
            I => \QuadInstance1.Quad_RNISL0OZ0Z_5\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__23511\,
            I => \N__23508\
        );

    \I__4254\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23505\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__23505\,
            I => \QuadInstance1.delayedCh_AZ0Z_2\
        );

    \I__4252\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23496\
        );

    \I__4251\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23496\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__23496\,
            I => \QuadInstance1.delayedCh_BZ0Z_2\
        );

    \I__4249\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23484\
        );

    \I__4248\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23484\
        );

    \I__4247\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23484\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__23484\,
            I => \QuadInstance1.delayedCh_AZ0Z_1\
        );

    \I__4245\ : CascadeMux
    port map (
            O => \N__23481\,
            I => \N__23478\
        );

    \I__4244\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23475\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__23475\,
            I => \QuadInstance1.Quad_RNI0Q0OZ0Z_9\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__23472\,
            I => \N__23469\
        );

    \I__4241\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23466\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__23466\,
            I => \QuadInstance1.Quad_RNI8P5DZ0Z_10\
        );

    \I__4239\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23460\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23455\
        );

    \I__4237\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23452\
        );

    \I__4236\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23445\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__23455\,
            I => \N__23441\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__23452\,
            I => \N__23438\
        );

    \I__4233\ : InMux
    port map (
            O => \N__23451\,
            I => \N__23435\
        );

    \I__4232\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23430\
        );

    \I__4231\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23430\
        );

    \I__4230\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23425\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__23445\,
            I => \N__23422\
        );

    \I__4228\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23419\
        );

    \I__4227\ : Span4Mux_h
    port map (
            O => \N__23441\,
            I => \N__23410\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__23438\,
            I => \N__23410\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__23435\,
            I => \N__23410\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__23430\,
            I => \N__23410\
        );

    \I__4223\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23405\
        );

    \I__4222\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23405\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__23425\,
            I => \N__23402\
        );

    \I__4220\ : Span4Mux_h
    port map (
            O => \N__23422\,
            I => \N__23397\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23397\
        );

    \I__4218\ : Span4Mux_v
    port map (
            O => \N__23410\,
            I => \N__23392\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__23405\,
            I => \N__23392\
        );

    \I__4216\ : Span4Mux_v
    port map (
            O => \N__23402\,
            I => \N__23388\
        );

    \I__4215\ : Span4Mux_v
    port map (
            O => \N__23397\,
            I => \N__23385\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__23392\,
            I => \N__23382\
        );

    \I__4213\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23379\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__23388\,
            I => \data_received_esr_RNIMIH31Z0Z_19\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__23385\,
            I => \data_received_esr_RNIMIH31Z0Z_19\
        );

    \I__4210\ : Odrv4
    port map (
            O => \N__23382\,
            I => \data_received_esr_RNIMIH31Z0Z_19\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__23379\,
            I => \data_received_esr_RNIMIH31Z0Z_19\
        );

    \I__4208\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23367\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__23367\,
            I => \N__23363\
        );

    \I__4206\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23359\
        );

    \I__4205\ : Span4Mux_v
    port map (
            O => \N__23363\,
            I => \N__23356\
        );

    \I__4204\ : InMux
    port map (
            O => \N__23362\,
            I => \N__23353\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__23359\,
            I => \N__23350\
        );

    \I__4202\ : Span4Mux_v
    port map (
            O => \N__23356\,
            I => \N__23345\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__23353\,
            I => \N__23345\
        );

    \I__4200\ : Odrv12
    port map (
            O => \N__23350\,
            I => \dataRead1_11\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__23345\,
            I => \dataRead1_11\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__23340\,
            I => \N__23337\
        );

    \I__4197\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23334\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__23334\,
            I => \QuadInstance1.Quad_RNI9Q5DZ0Z_11\
        );

    \I__4195\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23328\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__23328\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_11\
        );

    \I__4193\ : InMux
    port map (
            O => \N__23325\,
            I => \N__23322\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__23322\,
            I => \N__23319\
        );

    \I__4191\ : Span4Mux_h
    port map (
            O => \N__23319\,
            I => \N__23316\
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__23316\,
            I => \ch2_B_c\
        );

    \I__4189\ : InMux
    port map (
            O => \N__23313\,
            I => \N__23310\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__23310\,
            I => \N__23307\
        );

    \I__4187\ : Span4Mux_h
    port map (
            O => \N__23307\,
            I => \N__23304\
        );

    \I__4186\ : Sp12to4
    port map (
            O => \N__23304\,
            I => \N__23301\
        );

    \I__4185\ : Span12Mux_v
    port map (
            O => \N__23301\,
            I => \N__23298\
        );

    \I__4184\ : Odrv12
    port map (
            O => \N__23298\,
            I => \QuadInstance2.delayedCh_BZ0Z_0\
        );

    \I__4183\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23292\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__23292\,
            I => \N__23289\
        );

    \I__4181\ : Span4Mux_h
    port map (
            O => \N__23289\,
            I => \N__23286\
        );

    \I__4180\ : Span4Mux_h
    port map (
            O => \N__23286\,
            I => \N__23283\
        );

    \I__4179\ : Odrv4
    port map (
            O => \N__23283\,
            I => \ch4_B_c\
        );

    \I__4178\ : InMux
    port map (
            O => \N__23280\,
            I => \N__23277\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__23277\,
            I => \N__23274\
        );

    \I__4176\ : Span4Mux_h
    port map (
            O => \N__23274\,
            I => \N__23271\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__23271\,
            I => \N__23268\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__23268\,
            I => \ch4_A_c\
        );

    \I__4173\ : CascadeMux
    port map (
            O => \N__23265\,
            I => \N__23260\
        );

    \I__4172\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23257\
        );

    \I__4171\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23254\
        );

    \I__4170\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23251\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__23257\,
            I => \N__23246\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__23254\,
            I => \N__23246\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__23251\,
            I => \dataRead1_4\
        );

    \I__4166\ : Odrv4
    port map (
            O => \N__23246\,
            I => \dataRead1_4\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__23241\,
            I => \N__23238\
        );

    \I__4164\ : InMux
    port map (
            O => \N__23238\,
            I => \N__23235\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__23235\,
            I => \QuadInstance1.Quad_RNIRK0OZ0Z_4\
        );

    \I__4162\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23228\
        );

    \I__4161\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23225\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__23228\,
            I => \N__23222\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__23225\,
            I => \QuadInstance1.delayedCh_BZ0Z_1\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__23222\,
            I => \QuadInstance1.delayedCh_BZ0Z_1\
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__23217\,
            I => \PWMInstance4.un1_periodCounter12_1_0_a2_0_0_cascade_\
        );

    \I__4156\ : InMux
    port map (
            O => \N__23214\,
            I => \N__23211\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__23211\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_4\
        );

    \I__4154\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23205\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__23205\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_5\
        );

    \I__4152\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23199\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__23199\,
            I => \PWMInstance4.PWMPulseWidthCountZ0Z_10\
        );

    \I__4150\ : InMux
    port map (
            O => \N__23196\,
            I => \N__23192\
        );

    \I__4149\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23189\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__23192\,
            I => \N__23183\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__23189\,
            I => \N__23183\
        );

    \I__4146\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23180\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__23183\,
            I => \PWMInstance6.periodCounterZ0Z_15\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__23180\,
            I => \PWMInstance6.periodCounterZ0Z_15\
        );

    \I__4143\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23171\
        );

    \I__4142\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23168\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__23171\,
            I => \N__23162\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23162\
        );

    \I__4139\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23159\
        );

    \I__4138\ : Odrv4
    port map (
            O => \N__23162\,
            I => \PWMInstance6.periodCounterZ0Z_14\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__23159\,
            I => \PWMInstance6.periodCounterZ0Z_14\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__23154\,
            I => \N__23151\
        );

    \I__4135\ : InMux
    port map (
            O => \N__23151\,
            I => \N__23148\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__23148\,
            I => \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_5\
        );

    \I__4133\ : InMux
    port map (
            O => \N__23145\,
            I => \N__23142\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__23142\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_14\
        );

    \I__4131\ : CascadeMux
    port map (
            O => \N__23139\,
            I => \N__23136\
        );

    \I__4130\ : InMux
    port map (
            O => \N__23136\,
            I => \N__23133\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__23133\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_15\
        );

    \I__4128\ : InMux
    port map (
            O => \N__23130\,
            I => \N__23125\
        );

    \I__4127\ : InMux
    port map (
            O => \N__23129\,
            I => \N__23122\
        );

    \I__4126\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23119\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__23125\,
            I => \N__23116\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__23122\,
            I => \PWMInstance6.periodCounterZ0Z_10\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__23119\,
            I => \PWMInstance6.periodCounterZ0Z_10\
        );

    \I__4122\ : Odrv12
    port map (
            O => \N__23116\,
            I => \PWMInstance6.periodCounterZ0Z_10\
        );

    \I__4121\ : InMux
    port map (
            O => \N__23109\,
            I => \N__23106\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__23106\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_11\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__23103\,
            I => \N__23099\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__23102\,
            I => \N__23095\
        );

    \I__4117\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23092\
        );

    \I__4116\ : InMux
    port map (
            O => \N__23098\,
            I => \N__23089\
        );

    \I__4115\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23086\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__23092\,
            I => \N__23083\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__23089\,
            I => \PWMInstance6.periodCounterZ0Z_11\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__23086\,
            I => \PWMInstance6.periodCounterZ0Z_11\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__23083\,
            I => \PWMInstance6.periodCounterZ0Z_11\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__23076\,
            I => \N__23073\
        );

    \I__4109\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23070\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__23070\,
            I => \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_5\
        );

    \I__4107\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23064\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__23064\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_10\
        );

    \I__4105\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__23058\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_13\
        );

    \I__4103\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23050\
        );

    \I__4102\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23047\
        );

    \I__4101\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23044\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__23050\,
            I => \N__23041\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__23047\,
            I => \PWMInstance6.periodCounterZ0Z_12\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__23044\,
            I => \PWMInstance6.periodCounterZ0Z_12\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__23041\,
            I => \PWMInstance6.periodCounterZ0Z_12\
        );

    \I__4096\ : CascadeMux
    port map (
            O => \N__23034\,
            I => \N__23031\
        );

    \I__4095\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23027\
        );

    \I__4094\ : InMux
    port map (
            O => \N__23030\,
            I => \N__23023\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__23027\,
            I => \N__23020\
        );

    \I__4092\ : InMux
    port map (
            O => \N__23026\,
            I => \N__23017\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__23023\,
            I => \PWMInstance6.periodCounterZ0Z_13\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__23020\,
            I => \PWMInstance6.periodCounterZ0Z_13\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__23017\,
            I => \PWMInstance6.periodCounterZ0Z_13\
        );

    \I__4088\ : InMux
    port map (
            O => \N__23010\,
            I => \N__23007\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__23007\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_12\
        );

    \I__4086\ : InMux
    port map (
            O => \N__23004\,
            I => \N__23001\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__23001\,
            I => \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_5\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__22998\,
            I => \data_received_esr_RNIMIH31Z0Z_19_cascade_\
        );

    \I__4083\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22990\
        );

    \I__4082\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22985\
        );

    \I__4081\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22985\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__22990\,
            I => \data_receivedZ0Z_19\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__22985\,
            I => \data_receivedZ0Z_19\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__22980\,
            I => \N__22975\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__22979\,
            I => \N__22972\
        );

    \I__4076\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22965\
        );

    \I__4075\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22965\
        );

    \I__4074\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22965\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__22965\,
            I => \data_receivedZ0Z_23\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__22962\,
            I => \data_received_esr_RNIMIH31_0Z0Z_19_cascade_\
        );

    \I__4071\ : InMux
    port map (
            O => \N__22959\,
            I => \N__22956\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__22956\,
            I => \N__22953\
        );

    \I__4069\ : Span4Mux_h
    port map (
            O => \N__22953\,
            I => \N__22950\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__22950\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_5\
        );

    \I__4067\ : InMux
    port map (
            O => \N__22947\,
            I => \N__22944\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__22944\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_8\
        );

    \I__4065\ : InMux
    port map (
            O => \N__22941\,
            I => \N__22938\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__22938\,
            I => \N__22935\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__22935\,
            I => \OutRegZ0Z_11\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__22932\,
            I => \OutReg_esr_RNO_0Z0Z_12_cascade_\
        );

    \I__4061\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22926\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__22926\,
            I => \OutRegZ0Z_12\
        );

    \I__4059\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22919\
        );

    \I__4058\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22916\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__22919\,
            I => \data_receivedZ0Z_12\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__22916\,
            I => \data_receivedZ0Z_12\
        );

    \I__4055\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22907\
        );

    \I__4054\ : InMux
    port map (
            O => \N__22910\,
            I => \N__22904\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__22907\,
            I => \data_receivedZ0Z_13\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__22904\,
            I => \data_receivedZ0Z_13\
        );

    \I__4051\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22895\
        );

    \I__4050\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22892\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__22895\,
            I => \data_receivedZ0Z_14\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__22892\,
            I => \data_receivedZ0Z_14\
        );

    \I__4047\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22883\
        );

    \I__4046\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22880\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__22883\,
            I => \data_receivedZ0Z_10\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__22880\,
            I => \data_receivedZ0Z_10\
        );

    \I__4043\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22871\
        );

    \I__4042\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22868\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__22871\,
            I => \data_receivedZ0Z_11\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__22868\,
            I => \data_receivedZ0Z_11\
        );

    \I__4039\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22858\
        );

    \I__4038\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22855\
        );

    \I__4037\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22852\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__22858\,
            I => \QuadInstance6.delayedCh_AZ0Z_1\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__22855\,
            I => \QuadInstance6.delayedCh_AZ0Z_1\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__22852\,
            I => \QuadInstance6.delayedCh_AZ0Z_1\
        );

    \I__4033\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__22842\,
            I => \QuadInstance6.delayedCh_AZ0Z_2\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__22839\,
            I => \N__22835\
        );

    \I__4030\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22832\
        );

    \I__4029\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22829\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__22832\,
            I => \N__22826\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__22829\,
            I => \N__22823\
        );

    \I__4026\ : Span4Mux_v
    port map (
            O => \N__22826\,
            I => \N__22819\
        );

    \I__4025\ : Span4Mux_h
    port map (
            O => \N__22823\,
            I => \N__22816\
        );

    \I__4024\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22813\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__22819\,
            I => \dataRead6_13\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__22816\,
            I => \dataRead6_13\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__22813\,
            I => \dataRead6_13\
        );

    \I__4020\ : InMux
    port map (
            O => \N__22806\,
            I => \N__22802\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__22805\,
            I => \N__22799\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22784\
        );

    \I__4017\ : InMux
    port map (
            O => \N__22799\,
            I => \N__22780\
        );

    \I__4016\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22777\
        );

    \I__4015\ : InMux
    port map (
            O => \N__22797\,
            I => \N__22772\
        );

    \I__4014\ : InMux
    port map (
            O => \N__22796\,
            I => \N__22772\
        );

    \I__4013\ : InMux
    port map (
            O => \N__22795\,
            I => \N__22765\
        );

    \I__4012\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22765\
        );

    \I__4011\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22765\
        );

    \I__4010\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22762\
        );

    \I__4009\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22759\
        );

    \I__4008\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22750\
        );

    \I__4007\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22743\
        );

    \I__4006\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22743\
        );

    \I__4005\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22743\
        );

    \I__4004\ : Span4Mux_v
    port map (
            O => \N__22784\,
            I => \N__22740\
        );

    \I__4003\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22737\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22730\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__22777\,
            I => \N__22730\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__22772\,
            I => \N__22730\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__22765\,
            I => \N__22723\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__22762\,
            I => \N__22723\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__22759\,
            I => \N__22723\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__22758\,
            I => \N__22714\
        );

    \I__3995\ : CascadeMux
    port map (
            O => \N__22757\,
            I => \N__22711\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__22756\,
            I => \N__22707\
        );

    \I__3993\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22701\
        );

    \I__3992\ : InMux
    port map (
            O => \N__22754\,
            I => \N__22698\
        );

    \I__3991\ : InMux
    port map (
            O => \N__22753\,
            I => \N__22695\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__22750\,
            I => \N__22688\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__22743\,
            I => \N__22688\
        );

    \I__3988\ : Span4Mux_h
    port map (
            O => \N__22740\,
            I => \N__22688\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__22737\,
            I => \N__22681\
        );

    \I__3986\ : Sp12to4
    port map (
            O => \N__22730\,
            I => \N__22681\
        );

    \I__3985\ : Span12Mux_s3_v
    port map (
            O => \N__22723\,
            I => \N__22681\
        );

    \I__3984\ : InMux
    port map (
            O => \N__22722\,
            I => \N__22676\
        );

    \I__3983\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22676\
        );

    \I__3982\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22667\
        );

    \I__3981\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22667\
        );

    \I__3980\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22667\
        );

    \I__3979\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22667\
        );

    \I__3978\ : InMux
    port map (
            O => \N__22714\,
            I => \N__22652\
        );

    \I__3977\ : InMux
    port map (
            O => \N__22711\,
            I => \N__22652\
        );

    \I__3976\ : InMux
    port map (
            O => \N__22710\,
            I => \N__22652\
        );

    \I__3975\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22652\
        );

    \I__3974\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22652\
        );

    \I__3973\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22652\
        );

    \I__3972\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22652\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__22701\,
            I => \quadWriteZ0Z_6\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__22698\,
            I => \quadWriteZ0Z_6\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__22695\,
            I => \quadWriteZ0Z_6\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__22688\,
            I => \quadWriteZ0Z_6\
        );

    \I__3967\ : Odrv12
    port map (
            O => \N__22681\,
            I => \quadWriteZ0Z_6\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__22676\,
            I => \quadWriteZ0Z_6\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__22667\,
            I => \quadWriteZ0Z_6\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__22652\,
            I => \quadWriteZ0Z_6\
        );

    \I__3963\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22627\
        );

    \I__3962\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22624\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__22633\,
            I => \N__22621\
        );

    \I__3960\ : CascadeMux
    port map (
            O => \N__22632\,
            I => \N__22618\
        );

    \I__3959\ : CascadeMux
    port map (
            O => \N__22631\,
            I => \N__22615\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__22630\,
            I => \N__22611\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N__22599\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__22624\,
            I => \N__22599\
        );

    \I__3955\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22594\
        );

    \I__3954\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22594\
        );

    \I__3953\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22587\
        );

    \I__3952\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22587\
        );

    \I__3951\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22587\
        );

    \I__3950\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22572\
        );

    \I__3949\ : InMux
    port map (
            O => \N__22609\,
            I => \N__22572\
        );

    \I__3948\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22572\
        );

    \I__3947\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22572\
        );

    \I__3946\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22572\
        );

    \I__3945\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22572\
        );

    \I__3944\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22572\
        );

    \I__3943\ : Odrv12
    port map (
            O => \N__22599\,
            I => \QuadInstance6.un1_count_enable_i_a2_0_1\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__22594\,
            I => \QuadInstance6.un1_count_enable_i_a2_0_1\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__22587\,
            I => \QuadInstance6.un1_count_enable_i_a2_0_1\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__22572\,
            I => \QuadInstance6.un1_count_enable_i_a2_0_1\
        );

    \I__3939\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22559\
        );

    \I__3938\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22556\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__22559\,
            I => \N__22543\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22543\
        );

    \I__3935\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22540\
        );

    \I__3934\ : CascadeMux
    port map (
            O => \N__22554\,
            I => \N__22535\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__22553\,
            I => \N__22530\
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__22552\,
            I => \N__22525\
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__22551\,
            I => \N__22522\
        );

    \I__3930\ : InMux
    port map (
            O => \N__22550\,
            I => \N__22519\
        );

    \I__3929\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22514\
        );

    \I__3928\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22514\
        );

    \I__3927\ : Span4Mux_s3_v
    port map (
            O => \N__22543\,
            I => \N__22509\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__22540\,
            I => \N__22509\
        );

    \I__3925\ : InMux
    port map (
            O => \N__22539\,
            I => \N__22500\
        );

    \I__3924\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22500\
        );

    \I__3923\ : InMux
    port map (
            O => \N__22535\,
            I => \N__22500\
        );

    \I__3922\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22500\
        );

    \I__3921\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22487\
        );

    \I__3920\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22487\
        );

    \I__3919\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22487\
        );

    \I__3918\ : InMux
    port map (
            O => \N__22528\,
            I => \N__22487\
        );

    \I__3917\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22487\
        );

    \I__3916\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22487\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__22519\,
            I => \QuadInstance6.count_enable\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__22514\,
            I => \QuadInstance6.count_enable\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__22509\,
            I => \QuadInstance6.count_enable\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__22500\,
            I => \QuadInstance6.count_enable\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__22487\,
            I => \QuadInstance6.count_enable\
        );

    \I__3910\ : InMux
    port map (
            O => \N__22476\,
            I => \N__22473\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__22473\,
            I => \N__22470\
        );

    \I__3908\ : Odrv4
    port map (
            O => \N__22470\,
            I => \QuadInstance6.Quad_RNIJHNB1Z0Z_13\
        );

    \I__3907\ : InMux
    port map (
            O => \N__22467\,
            I => \N__22463\
        );

    \I__3906\ : InMux
    port map (
            O => \N__22466\,
            I => \N__22460\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__22463\,
            I => \QuadInstance6.delayedCh_BZ0Z_1\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__22460\,
            I => \QuadInstance6.delayedCh_BZ0Z_1\
        );

    \I__3903\ : InMux
    port map (
            O => \N__22455\,
            I => \N__22452\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__22452\,
            I => \N__22447\
        );

    \I__3901\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22444\
        );

    \I__3900\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22441\
        );

    \I__3899\ : Span4Mux_v
    port map (
            O => \N__22447\,
            I => \N__22436\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__22444\,
            I => \N__22436\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__22441\,
            I => \N__22433\
        );

    \I__3896\ : Span4Mux_h
    port map (
            O => \N__22436\,
            I => \N__22430\
        );

    \I__3895\ : Span12Mux_h
    port map (
            O => \N__22433\,
            I => \N__22427\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__22430\,
            I => \dataRead2_11\
        );

    \I__3893\ : Odrv12
    port map (
            O => \N__22427\,
            I => \dataRead2_11\
        );

    \I__3892\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22419\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__22419\,
            I => \N__22415\
        );

    \I__3890\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22411\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__22415\,
            I => \N__22408\
        );

    \I__3888\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22405\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__22411\,
            I => \N__22402\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__22408\,
            I => \dataRead3_11\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__22405\,
            I => \dataRead3_11\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__22402\,
            I => \dataRead3_11\
        );

    \I__3883\ : InMux
    port map (
            O => \N__22395\,
            I => \N__22392\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__22392\,
            I => \OutReg_0_4_i_m3_i_m3_ns_1_11\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__22389\,
            I => \N__22386\
        );

    \I__3880\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22382\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__22385\,
            I => \N__22379\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22375\
        );

    \I__3877\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22372\
        );

    \I__3876\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22369\
        );

    \I__3875\ : Span4Mux_h
    port map (
            O => \N__22375\,
            I => \N__22366\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__22372\,
            I => \dataRead5_12\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__22369\,
            I => \dataRead5_12\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__22366\,
            I => \dataRead5_12\
        );

    \I__3871\ : InMux
    port map (
            O => \N__22359\,
            I => \N__22356\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__22356\,
            I => \N__22353\
        );

    \I__3869\ : Span4Mux_h
    port map (
            O => \N__22353\,
            I => \N__22348\
        );

    \I__3868\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22345\
        );

    \I__3867\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22342\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__22348\,
            I => \N__22339\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__22345\,
            I => \dataRead2_12\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__22342\,
            I => \dataRead2_12\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__22339\,
            I => \dataRead2_12\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__22332\,
            I => \N__22328\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__22331\,
            I => \N__22325\
        );

    \I__3860\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22322\
        );

    \I__3859\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22319\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22316\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22312\
        );

    \I__3856\ : Span4Mux_v
    port map (
            O => \N__22316\,
            I => \N__22309\
        );

    \I__3855\ : InMux
    port map (
            O => \N__22315\,
            I => \N__22306\
        );

    \I__3854\ : Span4Mux_h
    port map (
            O => \N__22312\,
            I => \N__22303\
        );

    \I__3853\ : Span4Mux_h
    port map (
            O => \N__22309\,
            I => \N__22298\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__22306\,
            I => \N__22298\
        );

    \I__3851\ : Odrv4
    port map (
            O => \N__22303\,
            I => \dataRead3_12\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__22298\,
            I => \dataRead3_12\
        );

    \I__3849\ : InMux
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__22290\,
            I => \N__22286\
        );

    \I__3847\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22283\
        );

    \I__3846\ : Span4Mux_h
    port map (
            O => \N__22286\,
            I => \N__22279\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__22283\,
            I => \N__22276\
        );

    \I__3844\ : InMux
    port map (
            O => \N__22282\,
            I => \N__22273\
        );

    \I__3843\ : Span4Mux_v
    port map (
            O => \N__22279\,
            I => \N__22268\
        );

    \I__3842\ : Span4Mux_h
    port map (
            O => \N__22276\,
            I => \N__22268\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__22273\,
            I => \dataRead6_12\
        );

    \I__3840\ : Odrv4
    port map (
            O => \N__22268\,
            I => \dataRead6_12\
        );

    \I__3839\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22259\
        );

    \I__3838\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22256\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__22259\,
            I => \N__22253\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__22256\,
            I => \N__22249\
        );

    \I__3835\ : Span4Mux_v
    port map (
            O => \N__22253\,
            I => \N__22246\
        );

    \I__3834\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22243\
        );

    \I__3833\ : Span4Mux_v
    port map (
            O => \N__22249\,
            I => \N__22236\
        );

    \I__3832\ : Span4Mux_h
    port map (
            O => \N__22246\,
            I => \N__22236\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__22243\,
            I => \N__22236\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__22236\,
            I => \dataRead7_12\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__22233\,
            I => \OutReg_0_4_i_m3_ns_1_12_cascade_\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__22230\,
            I => \OutReg_esr_RNO_1Z0Z_12_cascade_\
        );

    \I__3827\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22224\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__22224\,
            I => \OutReg_esr_RNO_2Z0Z_12\
        );

    \I__3825\ : InMux
    port map (
            O => \N__22221\,
            I => \N__22218\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__22218\,
            I => \N__22215\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__22215\,
            I => \N__22212\
        );

    \I__3822\ : Odrv4
    port map (
            O => \N__22212\,
            I => \QuadInstance6.Quad_RNO_0_6_9\
        );

    \I__3821\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22206\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__22206\,
            I => \N__22203\
        );

    \I__3819\ : Span4Mux_h
    port map (
            O => \N__22203\,
            I => \N__22200\
        );

    \I__3818\ : Span4Mux_h
    port map (
            O => \N__22200\,
            I => \N__22197\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__22197\,
            I => \QuadInstance2.Quad_RNO_0_1_1\
        );

    \I__3816\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22178\
        );

    \I__3815\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22178\
        );

    \I__3814\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22178\
        );

    \I__3813\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22175\
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__22190\,
            I => \N__22172\
        );

    \I__3811\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22168\
        );

    \I__3810\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22165\
        );

    \I__3809\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22160\
        );

    \I__3808\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22160\
        );

    \I__3807\ : InMux
    port map (
            O => \N__22185\,
            I => \N__22156\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__22178\,
            I => \N__22151\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__22175\,
            I => \N__22151\
        );

    \I__3804\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22147\
        );

    \I__3803\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22144\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__22168\,
            I => \N__22136\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__22165\,
            I => \N__22131\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__22160\,
            I => \N__22131\
        );

    \I__3799\ : InMux
    port map (
            O => \N__22159\,
            I => \N__22128\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__22156\,
            I => \N__22123\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__22151\,
            I => \N__22123\
        );

    \I__3796\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22120\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__22147\,
            I => \N__22117\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__22144\,
            I => \N__22114\
        );

    \I__3793\ : InMux
    port map (
            O => \N__22143\,
            I => \N__22111\
        );

    \I__3792\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22089\
        );

    \I__3791\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22089\
        );

    \I__3790\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22089\
        );

    \I__3789\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22089\
        );

    \I__3788\ : Span4Mux_h
    port map (
            O => \N__22136\,
            I => \N__22084\
        );

    \I__3787\ : Span4Mux_v
    port map (
            O => \N__22131\,
            I => \N__22084\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22077\
        );

    \I__3785\ : Span4Mux_h
    port map (
            O => \N__22123\,
            I => \N__22077\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__22120\,
            I => \N__22077\
        );

    \I__3783\ : Span4Mux_h
    port map (
            O => \N__22117\,
            I => \N__22070\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__22114\,
            I => \N__22070\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__22111\,
            I => \N__22070\
        );

    \I__3780\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22059\
        );

    \I__3779\ : InMux
    port map (
            O => \N__22109\,
            I => \N__22059\
        );

    \I__3778\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22059\
        );

    \I__3777\ : InMux
    port map (
            O => \N__22107\,
            I => \N__22059\
        );

    \I__3776\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22059\
        );

    \I__3775\ : InMux
    port map (
            O => \N__22105\,
            I => \N__22042\
        );

    \I__3774\ : InMux
    port map (
            O => \N__22104\,
            I => \N__22042\
        );

    \I__3773\ : InMux
    port map (
            O => \N__22103\,
            I => \N__22042\
        );

    \I__3772\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22042\
        );

    \I__3771\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22042\
        );

    \I__3770\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22042\
        );

    \I__3769\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22042\
        );

    \I__3768\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22042\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__22089\,
            I => \quadWriteZ0Z_2\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__22084\,
            I => \quadWriteZ0Z_2\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__22077\,
            I => \quadWriteZ0Z_2\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__22070\,
            I => \quadWriteZ0Z_2\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__22059\,
            I => \quadWriteZ0Z_2\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__22042\,
            I => \quadWriteZ0Z_2\
        );

    \I__3761\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22026\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__22026\,
            I => \N__22023\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__22023\,
            I => \QuadInstance3.Quad_RNO_0_2_1\
        );

    \I__3758\ : InMux
    port map (
            O => \N__22020\,
            I => \N__22009\
        );

    \I__3757\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22005\
        );

    \I__3756\ : InMux
    port map (
            O => \N__22018\,
            I => \N__21997\
        );

    \I__3755\ : InMux
    port map (
            O => \N__22017\,
            I => \N__21994\
        );

    \I__3754\ : InMux
    port map (
            O => \N__22016\,
            I => \N__21991\
        );

    \I__3753\ : InMux
    port map (
            O => \N__22015\,
            I => \N__21986\
        );

    \I__3752\ : InMux
    port map (
            O => \N__22014\,
            I => \N__21986\
        );

    \I__3751\ : InMux
    port map (
            O => \N__22013\,
            I => \N__21980\
        );

    \I__3750\ : InMux
    port map (
            O => \N__22012\,
            I => \N__21980\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__22009\,
            I => \N__21977\
        );

    \I__3748\ : InMux
    port map (
            O => \N__22008\,
            I => \N__21974\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__22005\,
            I => \N__21971\
        );

    \I__3746\ : InMux
    port map (
            O => \N__22004\,
            I => \N__21958\
        );

    \I__3745\ : InMux
    port map (
            O => \N__22003\,
            I => \N__21958\
        );

    \I__3744\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21958\
        );

    \I__3743\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21958\
        );

    \I__3742\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21958\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__21997\,
            I => \N__21949\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__21994\,
            I => \N__21949\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__21991\,
            I => \N__21949\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__21986\,
            I => \N__21949\
        );

    \I__3737\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21946\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21941\
        );

    \I__3735\ : Span4Mux_v
    port map (
            O => \N__21977\,
            I => \N__21941\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21936\
        );

    \I__3733\ : Span4Mux_h
    port map (
            O => \N__21971\,
            I => \N__21936\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__21970\,
            I => \N__21930\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__21969\,
            I => \N__21924\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__21958\,
            I => \N__21912\
        );

    \I__3729\ : Span4Mux_v
    port map (
            O => \N__21949\,
            I => \N__21912\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__21946\,
            I => \N__21905\
        );

    \I__3727\ : Span4Mux_h
    port map (
            O => \N__21941\,
            I => \N__21905\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__21936\,
            I => \N__21905\
        );

    \I__3725\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21900\
        );

    \I__3724\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21900\
        );

    \I__3723\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21897\
        );

    \I__3722\ : InMux
    port map (
            O => \N__21930\,
            I => \N__21894\
        );

    \I__3721\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21881\
        );

    \I__3720\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21881\
        );

    \I__3719\ : InMux
    port map (
            O => \N__21927\,
            I => \N__21881\
        );

    \I__3718\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21881\
        );

    \I__3717\ : InMux
    port map (
            O => \N__21923\,
            I => \N__21881\
        );

    \I__3716\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21881\
        );

    \I__3715\ : InMux
    port map (
            O => \N__21921\,
            I => \N__21870\
        );

    \I__3714\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21870\
        );

    \I__3713\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21870\
        );

    \I__3712\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21870\
        );

    \I__3711\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21870\
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__21912\,
            I => \quadWriteZ0Z_3\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__21905\,
            I => \quadWriteZ0Z_3\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__21900\,
            I => \quadWriteZ0Z_3\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__21897\,
            I => \quadWriteZ0Z_3\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__21894\,
            I => \quadWriteZ0Z_3\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__21881\,
            I => \quadWriteZ0Z_3\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__21870\,
            I => \quadWriteZ0Z_3\
        );

    \I__3703\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21852\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__3701\ : Odrv4
    port map (
            O => \N__21849\,
            I => \QuadInstance3.Quad_RNO_0_3_4\
        );

    \I__3700\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21842\
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__21845\,
            I => \N__21839\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__21842\,
            I => \N__21835\
        );

    \I__3697\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21832\
        );

    \I__3696\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21829\
        );

    \I__3695\ : Span4Mux_h
    port map (
            O => \N__21835\,
            I => \N__21826\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__21832\,
            I => \N__21823\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__21829\,
            I => \N__21820\
        );

    \I__3692\ : Odrv4
    port map (
            O => \N__21826\,
            I => \dataRead3_4\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__21823\,
            I => \dataRead3_4\
        );

    \I__3690\ : Odrv12
    port map (
            O => \N__21820\,
            I => \dataRead3_4\
        );

    \I__3689\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21810\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__21810\,
            I => \QuadInstance1.Quad_RNO_0_1_9\
        );

    \I__3687\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21804\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21796\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__21803\,
            I => \N__21788\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__21802\,
            I => \N__21783\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__21801\,
            I => \N__21778\
        );

    \I__3682\ : CascadeMux
    port map (
            O => \N__21800\,
            I => \N__21774\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__21799\,
            I => \N__21771\
        );

    \I__3680\ : Span12Mux_s8_v
    port map (
            O => \N__21796\,
            I => \N__21768\
        );

    \I__3679\ : InMux
    port map (
            O => \N__21795\,
            I => \N__21765\
        );

    \I__3678\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21758\
        );

    \I__3677\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21758\
        );

    \I__3676\ : InMux
    port map (
            O => \N__21792\,
            I => \N__21758\
        );

    \I__3675\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21755\
        );

    \I__3674\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21744\
        );

    \I__3673\ : InMux
    port map (
            O => \N__21787\,
            I => \N__21744\
        );

    \I__3672\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21744\
        );

    \I__3671\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21744\
        );

    \I__3670\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21744\
        );

    \I__3669\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21733\
        );

    \I__3668\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21733\
        );

    \I__3667\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21733\
        );

    \I__3666\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21733\
        );

    \I__3665\ : InMux
    port map (
            O => \N__21771\,
            I => \N__21733\
        );

    \I__3664\ : Odrv12
    port map (
            O => \N__21768\,
            I => \QuadInstance7.count_enable\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__21765\,
            I => \QuadInstance7.count_enable\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__21758\,
            I => \QuadInstance7.count_enable\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__21755\,
            I => \QuadInstance7.count_enable\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__21744\,
            I => \QuadInstance7.count_enable\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__21733\,
            I => \QuadInstance7.count_enable\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__21720\,
            I => \N__21716\
        );

    \I__3657\ : CascadeMux
    port map (
            O => \N__21719\,
            I => \N__21713\
        );

    \I__3656\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21710\
        );

    \I__3655\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21707\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__21710\,
            I => \QuadInstance6.delayedCh_BZ0Z_2\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__21707\,
            I => \QuadInstance6.delayedCh_BZ0Z_2\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__21702\,
            I => \N__21699\
        );

    \I__3651\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21696\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__21696\,
            I => \N__21693\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__21693\,
            I => \QuadInstance6.Quad_RNIGENB1Z0Z_10\
        );

    \I__3648\ : InMux
    port map (
            O => \N__21690\,
            I => \bfn_13_7_0_\
        );

    \I__3647\ : InMux
    port map (
            O => \N__21687\,
            I => \QuadInstance1.un1_Quad_cry_8\
        );

    \I__3646\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21681\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__21681\,
            I => \QuadInstance1.Quad_RNO_0_1_10\
        );

    \I__3644\ : InMux
    port map (
            O => \N__21678\,
            I => \QuadInstance1.un1_Quad_cry_9\
        );

    \I__3643\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21672\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__21672\,
            I => \N__21669\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__21669\,
            I => \QuadInstance1.Quad_RNO_0_1_11\
        );

    \I__3640\ : InMux
    port map (
            O => \N__21666\,
            I => \QuadInstance1.un1_Quad_cry_10\
        );

    \I__3639\ : InMux
    port map (
            O => \N__21663\,
            I => \QuadInstance1.un1_Quad_cry_11\
        );

    \I__3638\ : InMux
    port map (
            O => \N__21660\,
            I => \QuadInstance1.un1_Quad_cry_12\
        );

    \I__3637\ : InMux
    port map (
            O => \N__21657\,
            I => \N__21654\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__21654\,
            I => \QuadInstance1.Quad_RNO_0_1_14\
        );

    \I__3635\ : InMux
    port map (
            O => \N__21651\,
            I => \QuadInstance1.un1_Quad_cry_13\
        );

    \I__3634\ : InMux
    port map (
            O => \N__21648\,
            I => \QuadInstance1.un1_Quad_cry_14\
        );

    \I__3633\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21642\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__21642\,
            I => \N__21639\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__21639\,
            I => \QuadInstance1.Quad_RNO_0_0_1\
        );

    \I__3630\ : InMux
    port map (
            O => \N__21636\,
            I => \QuadInstance1.un1_Quad_cry_0\
        );

    \I__3629\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__21630\,
            I => \N__21627\
        );

    \I__3627\ : Span4Mux_h
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__3626\ : Span4Mux_h
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__21621\,
            I => \QuadInstance1.Quad_RNO_0_1_2\
        );

    \I__3624\ : InMux
    port map (
            O => \N__21618\,
            I => \QuadInstance1.un1_Quad_cry_1\
        );

    \I__3623\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21612\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__21612\,
            I => \N__21609\
        );

    \I__3621\ : Span4Mux_v
    port map (
            O => \N__21609\,
            I => \N__21606\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__21606\,
            I => \QuadInstance1.Quad_RNO_0_1_3\
        );

    \I__3619\ : InMux
    port map (
            O => \N__21603\,
            I => \QuadInstance1.un1_Quad_cry_2\
        );

    \I__3618\ : InMux
    port map (
            O => \N__21600\,
            I => \N__21597\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__21597\,
            I => \QuadInstance1.Quad_RNO_0_1_4\
        );

    \I__3616\ : InMux
    port map (
            O => \N__21594\,
            I => \QuadInstance1.un1_Quad_cry_3\
        );

    \I__3615\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21588\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__21588\,
            I => \N__21585\
        );

    \I__3613\ : Odrv4
    port map (
            O => \N__21585\,
            I => \QuadInstance1.Quad_RNO_0_1_5\
        );

    \I__3612\ : InMux
    port map (
            O => \N__21582\,
            I => \QuadInstance1.un1_Quad_cry_4\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__21579\,
            I => \N__21576\
        );

    \I__3610\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21573\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__21573\,
            I => \N__21570\
        );

    \I__3608\ : Odrv4
    port map (
            O => \N__21570\,
            I => \QuadInstance1.Quad_RNO_0_1_6\
        );

    \I__3607\ : InMux
    port map (
            O => \N__21567\,
            I => \QuadInstance1.un1_Quad_cry_5\
        );

    \I__3606\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21561\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21558\
        );

    \I__3604\ : Odrv4
    port map (
            O => \N__21558\,
            I => \QuadInstance1.Quad_RNO_0_1_7\
        );

    \I__3603\ : InMux
    port map (
            O => \N__21555\,
            I => \QuadInstance1.un1_Quad_cry_6\
        );

    \I__3602\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21549\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__21549\,
            I => \N__21546\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__21546\,
            I => \N__21543\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__21543\,
            I => \QuadInstance1.Quad_RNO_0_1_8\
        );

    \I__3598\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21537\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__21537\,
            I => \N__21534\
        );

    \I__3596\ : Span4Mux_v
    port map (
            O => \N__21534\,
            I => \N__21531\
        );

    \I__3595\ : Span4Mux_h
    port map (
            O => \N__21531\,
            I => \N__21528\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__21528\,
            I => \ch0_A_c\
        );

    \I__3593\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21522\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__21522\,
            I => \N__21519\
        );

    \I__3591\ : Span4Mux_h
    port map (
            O => \N__21519\,
            I => \N__21516\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__21516\,
            I => \QuadInstance3.Quad_RNO_0_3_6\
        );

    \I__3589\ : CascadeMux
    port map (
            O => \N__21513\,
            I => \N__21510\
        );

    \I__3588\ : InMux
    port map (
            O => \N__21510\,
            I => \N__21507\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__21507\,
            I => \QuadInstance6.Quad_RNO_0_6_4\
        );

    \I__3586\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21501\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__21501\,
            I => \N__21497\
        );

    \I__3584\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21493\
        );

    \I__3583\ : Span12Mux_v
    port map (
            O => \N__21497\,
            I => \N__21490\
        );

    \I__3582\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21487\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__21493\,
            I => \N__21484\
        );

    \I__3580\ : Odrv12
    port map (
            O => \N__21490\,
            I => \dataRead6_4\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__21487\,
            I => \dataRead6_4\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__21484\,
            I => \dataRead6_4\
        );

    \I__3577\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21474\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__21474\,
            I => \N__21471\
        );

    \I__3575\ : Span4Mux_v
    port map (
            O => \N__21471\,
            I => \N__21468\
        );

    \I__3574\ : Odrv4
    port map (
            O => \N__21468\,
            I => \QuadInstance7.Quad_RNO_0_7_4\
        );

    \I__3573\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21461\
        );

    \I__3572\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21458\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__21461\,
            I => \N__21455\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__21458\,
            I => \N__21452\
        );

    \I__3569\ : Span4Mux_v
    port map (
            O => \N__21455\,
            I => \N__21446\
        );

    \I__3568\ : Span4Mux_v
    port map (
            O => \N__21452\,
            I => \N__21446\
        );

    \I__3567\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21443\
        );

    \I__3566\ : Span4Mux_h
    port map (
            O => \N__21446\,
            I => \N__21440\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__21443\,
            I => \dataRead7_4\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__21440\,
            I => \dataRead7_4\
        );

    \I__3563\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21432\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__21432\,
            I => \N__21429\
        );

    \I__3561\ : Odrv12
    port map (
            O => \N__21429\,
            I => \PWMInstance6.un1_periodCounter12_1_0_a2_0\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__21426\,
            I => \N__21423\
        );

    \I__3559\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21417\
        );

    \I__3558\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21414\
        );

    \I__3557\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21407\
        );

    \I__3556\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21407\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__21417\,
            I => \N__21404\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__21414\,
            I => \N__21401\
        );

    \I__3553\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21398\
        );

    \I__3552\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21395\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__21407\,
            I => \N__21390\
        );

    \I__3550\ : Span4Mux_v
    port map (
            O => \N__21404\,
            I => \N__21390\
        );

    \I__3549\ : Odrv4
    port map (
            O => \N__21401\,
            I => \PWMInstance6.out_0_sqmuxa\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__21398\,
            I => \PWMInstance6.out_0_sqmuxa\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__21395\,
            I => \PWMInstance6.out_0_sqmuxa\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__21390\,
            I => \PWMInstance6.out_0_sqmuxa\
        );

    \I__3545\ : InMux
    port map (
            O => \N__21381\,
            I => \bfn_12_17_0_\
        );

    \I__3544\ : IoInMux
    port map (
            O => \N__21378\,
            I => \N__21375\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__21375\,
            I => \N__21372\
        );

    \I__3542\ : Span4Mux_s1_v
    port map (
            O => \N__21372\,
            I => \N__21369\
        );

    \I__3541\ : Span4Mux_h
    port map (
            O => \N__21369\,
            I => \N__21365\
        );

    \I__3540\ : InMux
    port map (
            O => \N__21368\,
            I => \N__21362\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__21365\,
            I => \PWM6_c\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__21362\,
            I => \PWM6_c\
        );

    \I__3537\ : IoInMux
    port map (
            O => \N__21357\,
            I => \N__21354\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__21354\,
            I => \PWM5_obufLegalizeSB_DFFNet\
        );

    \I__3535\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21348\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__21348\,
            I => \N__21345\
        );

    \I__3533\ : Span4Mux_h
    port map (
            O => \N__21345\,
            I => \N__21342\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__21342\,
            I => \ch2_A_c\
        );

    \I__3531\ : InMux
    port map (
            O => \N__21339\,
            I => \N__21336\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__21336\,
            I => \N__21333\
        );

    \I__3529\ : Span12Mux_h
    port map (
            O => \N__21333\,
            I => \N__21330\
        );

    \I__3528\ : Odrv12
    port map (
            O => \N__21330\,
            I => \QuadInstance2.delayedCh_AZ0Z_0\
        );

    \I__3527\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21323\
        );

    \I__3526\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21320\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__21323\,
            I => \N__21317\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__21320\,
            I => \N__21313\
        );

    \I__3523\ : Span4Mux_v
    port map (
            O => \N__21317\,
            I => \N__21310\
        );

    \I__3522\ : InMux
    port map (
            O => \N__21316\,
            I => \N__21307\
        );

    \I__3521\ : Odrv12
    port map (
            O => \N__21313\,
            I => \dataRead5_4\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__21310\,
            I => \dataRead5_4\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__21307\,
            I => \dataRead5_4\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__21300\,
            I => \OutReg_ess_RNO_2Z0Z_4_cascade_\
        );

    \I__3517\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21292\
        );

    \I__3516\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21289\
        );

    \I__3515\ : InMux
    port map (
            O => \N__21295\,
            I => \N__21286\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__21292\,
            I => \N__21283\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__21289\,
            I => \N__21280\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__21286\,
            I => \N__21277\
        );

    \I__3511\ : Span12Mux_s9_h
    port map (
            O => \N__21283\,
            I => \N__21274\
        );

    \I__3510\ : Span4Mux_h
    port map (
            O => \N__21280\,
            I => \N__21271\
        );

    \I__3509\ : Span4Mux_v
    port map (
            O => \N__21277\,
            I => \N__21268\
        );

    \I__3508\ : Odrv12
    port map (
            O => \N__21274\,
            I => \dataRead2_4\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__21271\,
            I => \dataRead2_4\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__21268\,
            I => \dataRead2_4\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__21261\,
            I => \OutReg_0_4_i_m3_ns_1_4_cascade_\
        );

    \I__3504\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21255\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__21255\,
            I => \OutReg_ess_RNO_1Z0Z_4\
        );

    \I__3502\ : InMux
    port map (
            O => \N__21252\,
            I => \N__21249\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__21249\,
            I => \OutReg_0_5_i_m3_ns_1_4\
        );

    \I__3500\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21241\
        );

    \I__3499\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21238\
        );

    \I__3498\ : InMux
    port map (
            O => \N__21244\,
            I => \N__21235\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__21241\,
            I => \PWMInstance6.periodCounterZ0Z_8\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__21238\,
            I => \PWMInstance6.periodCounterZ0Z_8\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__21235\,
            I => \PWMInstance6.periodCounterZ0Z_8\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__21228\,
            I => \N__21223\
        );

    \I__3493\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21220\
        );

    \I__3492\ : InMux
    port map (
            O => \N__21226\,
            I => \N__21217\
        );

    \I__3491\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21214\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__21220\,
            I => \PWMInstance6.periodCounterZ0Z_9\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__21217\,
            I => \PWMInstance6.periodCounterZ0Z_9\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__21214\,
            I => \PWMInstance6.periodCounterZ0Z_9\
        );

    \I__3487\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21204\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__21204\,
            I => \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_5\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__21201\,
            I => \N__21198\
        );

    \I__3484\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21195\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__21195\,
            I => \N__21192\
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__21192\,
            I => \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_5\
        );

    \I__3481\ : InMux
    port map (
            O => \N__21189\,
            I => \N__21186\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21183\
        );

    \I__3479\ : Odrv4
    port map (
            O => \N__21183\,
            I => \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_5\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__21180\,
            I => \N__21177\
        );

    \I__3477\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21174\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__21174\,
            I => \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_5\
        );

    \I__3475\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21168\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__21168\,
            I => \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_5\
        );

    \I__3473\ : CascadeMux
    port map (
            O => \N__21165\,
            I => \PWMInstance6.un1_periodCounter12_1_0_a2_0_6_cascade_\
        );

    \I__3472\ : CascadeMux
    port map (
            O => \N__21162\,
            I => \N__21159\
        );

    \I__3471\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21155\
        );

    \I__3470\ : InMux
    port map (
            O => \N__21158\,
            I => \N__21151\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__21155\,
            I => \N__21148\
        );

    \I__3468\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21145\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__21151\,
            I => \PWMInstance6.periodCounter12\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__21148\,
            I => \PWMInstance6.periodCounter12\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__21145\,
            I => \PWMInstance6.periodCounter12\
        );

    \I__3464\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21135\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__21132\,
            I => \N__21129\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__21129\,
            I => \PWMInstance6.un1_periodCounter12_1_0_a2_0_14\
        );

    \I__3460\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21123\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__21123\,
            I => \N__21120\
        );

    \I__3458\ : Span4Mux_v
    port map (
            O => \N__21120\,
            I => \N__21117\
        );

    \I__3457\ : IoSpan4Mux
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__21114\,
            I => \ch6_A_c\
        );

    \I__3455\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21108\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__21108\,
            I => \N__21105\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__21105\,
            I => \N__21102\
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__21102\,
            I => \QuadInstance6.delayedCh_AZ0Z_0\
        );

    \I__3451\ : InMux
    port map (
            O => \N__21099\,
            I => \N__21096\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__21096\,
            I => \N__21093\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__21093\,
            I => \PWMInstance6.un1_periodCounter12_1_0_a2_0_9\
        );

    \I__3448\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21085\
        );

    \I__3447\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21080\
        );

    \I__3446\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21080\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__21085\,
            I => \PWMInstance6.periodCounterZ0Z_0\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__21080\,
            I => \PWMInstance6.periodCounterZ0Z_0\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__21075\,
            I => \N__21070\
        );

    \I__3442\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21067\
        );

    \I__3441\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21064\
        );

    \I__3440\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21061\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__21067\,
            I => \PWMInstance6.periodCounterZ0Z_1\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__21064\,
            I => \PWMInstance6.periodCounterZ0Z_1\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__21061\,
            I => \PWMInstance6.periodCounterZ0Z_1\
        );

    \I__3436\ : InMux
    port map (
            O => \N__21054\,
            I => \N__21051\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__21051\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_0\
        );

    \I__3434\ : InMux
    port map (
            O => \N__21048\,
            I => \N__21045\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__21045\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_1\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__21042\,
            I => \N__21038\
        );

    \I__3431\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21034\
        );

    \I__3430\ : InMux
    port map (
            O => \N__21038\,
            I => \N__21029\
        );

    \I__3429\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21029\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__21034\,
            I => \PWMInstance6.periodCounterZ0Z_6\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__21029\,
            I => \PWMInstance6.periodCounterZ0Z_6\
        );

    \I__3426\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21019\
        );

    \I__3425\ : InMux
    port map (
            O => \N__21023\,
            I => \N__21016\
        );

    \I__3424\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21013\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__21019\,
            I => \PWMInstance6.periodCounterZ0Z_7\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__21016\,
            I => \PWMInstance6.periodCounterZ0Z_7\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__21013\,
            I => \PWMInstance6.periodCounterZ0Z_7\
        );

    \I__3420\ : InMux
    port map (
            O => \N__21006\,
            I => \N__21003\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__21003\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_6\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__21000\,
            I => \N__20997\
        );

    \I__3417\ : InMux
    port map (
            O => \N__20997\,
            I => \N__20994\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__20994\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_7\
        );

    \I__3415\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20983\
        );

    \I__3414\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20983\
        );

    \I__3413\ : InMux
    port map (
            O => \N__20989\,
            I => \N__20978\
        );

    \I__3412\ : InMux
    port map (
            O => \N__20988\,
            I => \N__20978\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__20983\,
            I => \PWMInstance6.clkCountZ0Z_0\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__20978\,
            I => \PWMInstance6.clkCountZ0Z_0\
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__20973\,
            I => \N__20970\
        );

    \I__3408\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20962\
        );

    \I__3407\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20962\
        );

    \I__3406\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20957\
        );

    \I__3405\ : InMux
    port map (
            O => \N__20967\,
            I => \N__20957\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__20962\,
            I => \PWMInstance6.clkCountZ0Z_1\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__20957\,
            I => \PWMInstance6.clkCountZ0Z_1\
        );

    \I__3402\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20946\
        );

    \I__3401\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20946\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__20946\,
            I => \pwmWrite_fastZ0Z_6\
        );

    \I__3399\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20936\
        );

    \I__3398\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20936\
        );

    \I__3397\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20933\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__20936\,
            I => \pwmWriteZ0Z_6\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__20933\,
            I => \pwmWriteZ0Z_6\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__20928\,
            I => \N__20925\
        );

    \I__3393\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20918\
        );

    \I__3392\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20918\
        );

    \I__3391\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20915\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__20918\,
            I => \N__20912\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__20915\,
            I => \PWMInstance6.periodCounterZ0Z_16\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__20912\,
            I => \PWMInstance6.periodCounterZ0Z_16\
        );

    \I__3387\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__20904\,
            I => \data_receivedZ0Z_18\
        );

    \I__3385\ : InMux
    port map (
            O => \N__20901\,
            I => \N__20898\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__20898\,
            I => \data_receivedZ0Z_17\
        );

    \I__3383\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20892\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__20892\,
            I => \data_receivedZ0Z_16\
        );

    \I__3381\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20885\
        );

    \I__3380\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20882\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__20885\,
            I => \data_receivedZ0Z_15\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__20882\,
            I => \data_receivedZ0Z_15\
        );

    \I__3377\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20872\
        );

    \I__3376\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20869\
        );

    \I__3375\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20866\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__20872\,
            I => \N__20863\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__20869\,
            I => \N__20860\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20857\
        );

    \I__3371\ : Span4Mux_h
    port map (
            O => \N__20863\,
            I => \N__20852\
        );

    \I__3370\ : Span4Mux_h
    port map (
            O => \N__20860\,
            I => \N__20852\
        );

    \I__3369\ : Span4Mux_v
    port map (
            O => \N__20857\,
            I => \N__20849\
        );

    \I__3368\ : Odrv4
    port map (
            O => \N__20852\,
            I => \dataRead7_11\
        );

    \I__3367\ : Odrv4
    port map (
            O => \N__20849\,
            I => \dataRead7_11\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__20844\,
            I => \N__20841\
        );

    \I__3365\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20837\
        );

    \I__3364\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20834\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__20837\,
            I => \N__20831\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__20834\,
            I => \N__20825\
        );

    \I__3361\ : Span4Mux_v
    port map (
            O => \N__20831\,
            I => \N__20825\
        );

    \I__3360\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20822\
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__20825\,
            I => \dataRead6_11\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__20822\,
            I => \dataRead6_11\
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__20817\,
            I => \OutReg_ess_RNO_1Z0Z_11_cascade_\
        );

    \I__3356\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__20811\,
            I => \OutReg_ess_RNO_2Z0Z_11\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__20808\,
            I => \OutReg_ess_RNO_0Z0Z_11_cascade_\
        );

    \I__3353\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__20802\,
            I => \OutReg_ess_RNO_0Z0Z_13\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__3350\ : InMux
    port map (
            O => \N__20796\,
            I => \N__20793\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__20793\,
            I => \N__20790\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__20790\,
            I => \QuadInstance6.Quad_RNI79A91Z0Z_8\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__20787\,
            I => \QuadInstance6.un1_count_enable_i_a2_0_1_cascade_\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__20784\,
            I => \N__20781\
        );

    \I__3345\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20778\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__20778\,
            I => \N__20775\
        );

    \I__3343\ : Odrv12
    port map (
            O => \N__20775\,
            I => \QuadInstance6.Quad_RNI35A91Z0Z_4\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__20772\,
            I => \N__20769\
        );

    \I__3341\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20766\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__20766\,
            I => \N__20763\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__20763\,
            I => \QuadInstance6.Quad_RNIIGNB1Z0Z_12\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__20760\,
            I => \N__20757\
        );

    \I__3337\ : InMux
    port map (
            O => \N__20757\,
            I => \N__20754\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__20754\,
            I => \N__20751\
        );

    \I__3335\ : Odrv12
    port map (
            O => \N__20751\,
            I => \QuadInstance6.Quad_RNI57A91Z0Z_6\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__20748\,
            I => \N__20745\
        );

    \I__3333\ : InMux
    port map (
            O => \N__20745\,
            I => \N__20742\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__20742\,
            I => \N__20739\
        );

    \I__3331\ : Odrv12
    port map (
            O => \N__20739\,
            I => \QuadInstance6.Quad_RNI68A91Z0Z_7\
        );

    \I__3330\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20733\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__20733\,
            I => \OutReg_0_4_i_m3_ns_1_13\
        );

    \I__3328\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__20727\,
            I => \OutReg_ess_RNO_1Z0Z_13\
        );

    \I__3326\ : InMux
    port map (
            O => \N__20724\,
            I => \N__20721\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__20721\,
            I => \N__20718\
        );

    \I__3324\ : Span4Mux_v
    port map (
            O => \N__20718\,
            I => \N__20715\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__20715\,
            I => \QuadInstance7.Quad_RNO_0_7_10\
        );

    \I__3322\ : InMux
    port map (
            O => \N__20712\,
            I => \N__20709\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__20709\,
            I => \N__20706\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__20706\,
            I => \QuadInstance5.Quad_RNO_0_5_9\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__20703\,
            I => \N__20700\
        );

    \I__3318\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20697\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__20697\,
            I => \N__20694\
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__20694\,
            I => \QuadInstance6.Quad_RNI02A91Z0Z_1\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__20691\,
            I => \QuadInstance6.count_enable_cascade_\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__20688\,
            I => \N__20685\
        );

    \I__3313\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20682\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__20682\,
            I => \N__20679\
        );

    \I__3311\ : Odrv4
    port map (
            O => \N__20679\,
            I => \QuadInstance6.Quad_RNI13A91Z0Z_2\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__20676\,
            I => \N__20673\
        );

    \I__3309\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20670\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__20670\,
            I => \N__20667\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__20667\,
            I => \QuadInstance6.Quad_RNIHFNB1Z0Z_11\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__20664\,
            I => \N__20661\
        );

    \I__3305\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20658\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20655\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__20655\,
            I => \QuadInstance6.Quad_RNI24A91Z0Z_3\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__20652\,
            I => \N__20649\
        );

    \I__3301\ : InMux
    port map (
            O => \N__20649\,
            I => \N__20646\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__20646\,
            I => \N__20643\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__20643\,
            I => \QuadInstance6.Quad_RNI46A91Z0Z_5\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__20640\,
            I => \N__20637\
        );

    \I__3297\ : InMux
    port map (
            O => \N__20637\,
            I => \N__20634\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__20634\,
            I => \N__20631\
        );

    \I__3295\ : Odrv4
    port map (
            O => \N__20631\,
            I => \QuadInstance6.Quad_RNI8AA91Z0Z_9\
        );

    \I__3294\ : InMux
    port map (
            O => \N__20628\,
            I => \QuadInstance6.un1_Quad_cry_11\
        );

    \I__3293\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20622\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__20622\,
            I => \N__20619\
        );

    \I__3291\ : Odrv4
    port map (
            O => \N__20619\,
            I => \QuadInstance6.Quad_RNO_0_6_13\
        );

    \I__3290\ : InMux
    port map (
            O => \N__20616\,
            I => \QuadInstance6.un1_Quad_cry_12\
        );

    \I__3289\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20610\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__20610\,
            I => \N__20607\
        );

    \I__3287\ : Odrv12
    port map (
            O => \N__20607\,
            I => \QuadInstance6.Quad_RNIKINB1Z0Z_14\
        );

    \I__3286\ : InMux
    port map (
            O => \N__20604\,
            I => \QuadInstance6.un1_Quad_cry_13\
        );

    \I__3285\ : InMux
    port map (
            O => \N__20601\,
            I => \N__20598\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__20598\,
            I => \N__20595\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__20595\,
            I => \QuadInstance6.un1_Quad_axb_15\
        );

    \I__3282\ : InMux
    port map (
            O => \N__20592\,
            I => \QuadInstance6.un1_Quad_cry_14\
        );

    \I__3281\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20586\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__20586\,
            I => \N__20583\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__20583\,
            I => \QuadInstance6.Quad_RNO_0_5_1\
        );

    \I__3278\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20574\
        );

    \I__3276\ : Span4Mux_h
    port map (
            O => \N__20574\,
            I => \N__20571\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__20571\,
            I => \QuadInstance7.Quad_RNO_0_7_8\
        );

    \I__3274\ : InMux
    port map (
            O => \N__20568\,
            I => \N__20565\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__20565\,
            I => \QuadInstance6.Quad_RNO_0_6_14\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__20562\,
            I => \N__20559\
        );

    \I__3271\ : InMux
    port map (
            O => \N__20559\,
            I => \N__20555\
        );

    \I__3270\ : InMux
    port map (
            O => \N__20558\,
            I => \N__20551\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__20555\,
            I => \N__20548\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__20554\,
            I => \N__20545\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20542\
        );

    \I__3266\ : Span12Mux_s5_v
    port map (
            O => \N__20548\,
            I => \N__20539\
        );

    \I__3265\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20536\
        );

    \I__3264\ : Span4Mux_h
    port map (
            O => \N__20542\,
            I => \N__20533\
        );

    \I__3263\ : Odrv12
    port map (
            O => \N__20539\,
            I => \dataRead6_14\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__20536\,
            I => \dataRead6_14\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__20533\,
            I => \dataRead6_14\
        );

    \I__3260\ : InMux
    port map (
            O => \N__20526\,
            I => \N__20523\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__20523\,
            I => \QuadInstance6.Quad_RNO_0_6_10\
        );

    \I__3258\ : InMux
    port map (
            O => \N__20520\,
            I => \QuadInstance6.un1_Quad_cry_3\
        );

    \I__3257\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20514\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__20514\,
            I => \QuadInstance6.Quad_RNO_0_6_5\
        );

    \I__3255\ : InMux
    port map (
            O => \N__20511\,
            I => \QuadInstance6.un1_Quad_cry_4\
        );

    \I__3254\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20505\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__20505\,
            I => \QuadInstance6.Quad_RNO_0_6_6\
        );

    \I__3252\ : InMux
    port map (
            O => \N__20502\,
            I => \QuadInstance6.un1_Quad_cry_5\
        );

    \I__3251\ : InMux
    port map (
            O => \N__20499\,
            I => \N__20496\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__20496\,
            I => \QuadInstance6.Quad_RNO_0_6_7\
        );

    \I__3249\ : InMux
    port map (
            O => \N__20493\,
            I => \QuadInstance6.un1_Quad_cry_6\
        );

    \I__3248\ : InMux
    port map (
            O => \N__20490\,
            I => \N__20487\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__20487\,
            I => \QuadInstance6.Quad_RNO_0_6_8\
        );

    \I__3246\ : InMux
    port map (
            O => \N__20484\,
            I => \bfn_12_6_0_\
        );

    \I__3245\ : InMux
    port map (
            O => \N__20481\,
            I => \QuadInstance6.un1_Quad_cry_8\
        );

    \I__3244\ : InMux
    port map (
            O => \N__20478\,
            I => \QuadInstance6.un1_Quad_cry_9\
        );

    \I__3243\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20472\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__20472\,
            I => \QuadInstance6.Quad_RNO_0_6_11\
        );

    \I__3241\ : InMux
    port map (
            O => \N__20469\,
            I => \QuadInstance6.un1_Quad_cry_10\
        );

    \I__3240\ : InMux
    port map (
            O => \N__20466\,
            I => \N__20463\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__20463\,
            I => \N__20460\
        );

    \I__3238\ : Odrv4
    port map (
            O => \N__20460\,
            I => \QuadInstance6.Quad_RNO_0_6_12\
        );

    \I__3237\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20454\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__20454\,
            I => \N__20451\
        );

    \I__3235\ : Span4Mux_h
    port map (
            O => \N__20451\,
            I => \N__20448\
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__20448\,
            I => \QuadInstance5.Quad_RNO_0_5_5\
        );

    \I__3233\ : InMux
    port map (
            O => \N__20445\,
            I => \N__20442\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__20442\,
            I => \N__20439\
        );

    \I__3231\ : Span4Mux_h
    port map (
            O => \N__20439\,
            I => \N__20436\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__20436\,
            I => \QuadInstance7.Quad_RNO_0_7_5\
        );

    \I__3229\ : InMux
    port map (
            O => \N__20433\,
            I => \QuadInstance6.un1_Quad_cry_0\
        );

    \I__3228\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20427\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__20427\,
            I => \QuadInstance6.Quad_RNO_0_6_2\
        );

    \I__3226\ : InMux
    port map (
            O => \N__20424\,
            I => \QuadInstance6.un1_Quad_cry_1\
        );

    \I__3225\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20418\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__20418\,
            I => \QuadInstance6.Quad_RNO_0_6_3\
        );

    \I__3223\ : InMux
    port map (
            O => \N__20415\,
            I => \QuadInstance6.un1_Quad_cry_2\
        );

    \I__3222\ : InMux
    port map (
            O => \N__20412\,
            I => \PWMInstance6.un1_periodCounter_2_cry_12\
        );

    \I__3221\ : InMux
    port map (
            O => \N__20409\,
            I => \PWMInstance6.un1_periodCounter_2_cry_13\
        );

    \I__3220\ : InMux
    port map (
            O => \N__20406\,
            I => \PWMInstance6.un1_periodCounter_2_cry_14\
        );

    \I__3219\ : InMux
    port map (
            O => \N__20403\,
            I => \bfn_11_16_0_\
        );

    \I__3218\ : InMux
    port map (
            O => \N__20400\,
            I => \N__20397\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__20397\,
            I => \N__20394\
        );

    \I__3216\ : Span4Mux_h
    port map (
            O => \N__20394\,
            I => \N__20391\
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__20391\,
            I => \ch3_A_c\
        );

    \I__3214\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20385\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__20385\,
            I => \N__20382\
        );

    \I__3212\ : Span4Mux_v
    port map (
            O => \N__20382\,
            I => \N__20379\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__20379\,
            I => \N__20376\
        );

    \I__3210\ : Span4Mux_v
    port map (
            O => \N__20376\,
            I => \N__20373\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__20373\,
            I => \QuadInstance3.delayedCh_AZ0Z_0\
        );

    \I__3208\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20367\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__20367\,
            I => \N__20364\
        );

    \I__3206\ : Span4Mux_h
    port map (
            O => \N__20364\,
            I => \N__20361\
        );

    \I__3205\ : Span4Mux_h
    port map (
            O => \N__20361\,
            I => \N__20358\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__20358\,
            I => \QuadInstance2.Quad_RNO_0_2_5\
        );

    \I__3203\ : InMux
    port map (
            O => \N__20355\,
            I => \N__20352\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__20352\,
            I => \N__20347\
        );

    \I__3201\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20344\
        );

    \I__3200\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20341\
        );

    \I__3199\ : Span4Mux_v
    port map (
            O => \N__20347\,
            I => \N__20338\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__20344\,
            I => \PWMInstance6.periodCounterZ0Z_4\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__20341\,
            I => \PWMInstance6.periodCounterZ0Z_4\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__20338\,
            I => \PWMInstance6.periodCounterZ0Z_4\
        );

    \I__3195\ : InMux
    port map (
            O => \N__20331\,
            I => \PWMInstance6.un1_periodCounter_2_cry_3\
        );

    \I__3194\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20324\
        );

    \I__3193\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20320\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__20324\,
            I => \N__20317\
        );

    \I__3191\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20314\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__20320\,
            I => \PWMInstance6.periodCounterZ0Z_5\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__20317\,
            I => \PWMInstance6.periodCounterZ0Z_5\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__20314\,
            I => \PWMInstance6.periodCounterZ0Z_5\
        );

    \I__3187\ : InMux
    port map (
            O => \N__20307\,
            I => \PWMInstance6.un1_periodCounter_2_cry_4\
        );

    \I__3186\ : InMux
    port map (
            O => \N__20304\,
            I => \PWMInstance6.un1_periodCounter_2_cry_5\
        );

    \I__3185\ : InMux
    port map (
            O => \N__20301\,
            I => \PWMInstance6.un1_periodCounter_2_cry_6\
        );

    \I__3184\ : InMux
    port map (
            O => \N__20298\,
            I => \bfn_11_15_0_\
        );

    \I__3183\ : InMux
    port map (
            O => \N__20295\,
            I => \PWMInstance6.un1_periodCounter_2_cry_8\
        );

    \I__3182\ : InMux
    port map (
            O => \N__20292\,
            I => \PWMInstance6.un1_periodCounter_2_cry_9\
        );

    \I__3181\ : InMux
    port map (
            O => \N__20289\,
            I => \PWMInstance6.un1_periodCounter_2_cry_10\
        );

    \I__3180\ : InMux
    port map (
            O => \N__20286\,
            I => \PWMInstance6.un1_periodCounter_2_cry_11\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__20283\,
            I => \N__20279\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__20282\,
            I => \N__20276\
        );

    \I__3177\ : InMux
    port map (
            O => \N__20279\,
            I => \N__20273\
        );

    \I__3176\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20270\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__20273\,
            I => \N__20267\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__20270\,
            I => \N__20264\
        );

    \I__3173\ : Span4Mux_v
    port map (
            O => \N__20267\,
            I => \N__20260\
        );

    \I__3172\ : Span4Mux_h
    port map (
            O => \N__20264\,
            I => \N__20257\
        );

    \I__3171\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20254\
        );

    \I__3170\ : Odrv4
    port map (
            O => \N__20260\,
            I => \dataRead7_14\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__20257\,
            I => \dataRead7_14\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__20254\,
            I => \dataRead7_14\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__20247\,
            I => \OutReg_0_4_i_m3_ns_1_14_cascade_\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__20244\,
            I => \N__20241\
        );

    \I__3165\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20235\
        );

    \I__3164\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20235\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__20235\,
            I => \pwmWrite_fastZ0Z_5\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__20232\,
            I => \N__20228\
        );

    \I__3161\ : CascadeMux
    port map (
            O => \N__20231\,
            I => \N__20225\
        );

    \I__3160\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20217\
        );

    \I__3159\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20217\
        );

    \I__3158\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20217\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__20217\,
            I => \pwmWriteZ0Z_5\
        );

    \I__3156\ : InMux
    port map (
            O => \N__20214\,
            I => \PWMInstance6.un1_periodCounter_2_cry_0\
        );

    \I__3155\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20206\
        );

    \I__3154\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20203\
        );

    \I__3153\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20200\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__20206\,
            I => \N__20197\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__20203\,
            I => \PWMInstance6.periodCounterZ0Z_2\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__20200\,
            I => \PWMInstance6.periodCounterZ0Z_2\
        );

    \I__3149\ : Odrv4
    port map (
            O => \N__20197\,
            I => \PWMInstance6.periodCounterZ0Z_2\
        );

    \I__3148\ : InMux
    port map (
            O => \N__20190\,
            I => \PWMInstance6.un1_periodCounter_2_cry_1\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__20187\,
            I => \N__20184\
        );

    \I__3146\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__20181\,
            I => \N__20176\
        );

    \I__3144\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20173\
        );

    \I__3143\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20170\
        );

    \I__3142\ : Span4Mux_v
    port map (
            O => \N__20176\,
            I => \N__20167\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__20173\,
            I => \PWMInstance6.periodCounterZ0Z_3\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__20170\,
            I => \PWMInstance6.periodCounterZ0Z_3\
        );

    \I__3139\ : Odrv4
    port map (
            O => \N__20167\,
            I => \PWMInstance6.periodCounterZ0Z_3\
        );

    \I__3138\ : InMux
    port map (
            O => \N__20160\,
            I => \PWMInstance6.un1_periodCounter_2_cry_2\
        );

    \I__3137\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20154\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__20154\,
            I => \QuadInstance3.Quad_RNO_0_3_14\
        );

    \I__3135\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20148\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__20148\,
            I => \N__20145\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__20145\,
            I => \QuadInstance5.Quad_RNO_0_5_2\
        );

    \I__3132\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20139\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__20139\,
            I => \N__20136\
        );

    \I__3130\ : Odrv4
    port map (
            O => \N__20136\,
            I => \QuadInstance7.Quad_RNO_0_7_14\
        );

    \I__3129\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20130\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__20130\,
            I => \QuadInstance3.Quad_RNO_0_3_10\
        );

    \I__3127\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20124\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__20124\,
            I => \QuadInstance3.Quad_RNO_0_3_11\
        );

    \I__3125\ : InMux
    port map (
            O => \N__20121\,
            I => \N__20118\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__20118\,
            I => \N__20115\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__20115\,
            I => \OutReg_ess_RNO_2Z0Z_13\
        );

    \I__3122\ : InMux
    port map (
            O => \N__20112\,
            I => \N__20109\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__20109\,
            I => \N__20105\
        );

    \I__3120\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20102\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__20105\,
            I => \N__20098\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__20102\,
            I => \N__20095\
        );

    \I__3117\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20092\
        );

    \I__3116\ : Span4Mux_h
    port map (
            O => \N__20098\,
            I => \N__20087\
        );

    \I__3115\ : Span4Mux_h
    port map (
            O => \N__20095\,
            I => \N__20087\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__20092\,
            I => \dataRead5_11\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__20087\,
            I => \dataRead5_11\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__20082\,
            I => \OutReg_0_5_i_m3_i_m3_ns_1_11_cascade_\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__20079\,
            I => \N__20076\
        );

    \I__3110\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20073\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__20073\,
            I => \N__20069\
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__20072\,
            I => \N__20066\
        );

    \I__3107\ : Span4Mux_v
    port map (
            O => \N__20069\,
            I => \N__20062\
        );

    \I__3106\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20059\
        );

    \I__3105\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20056\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__20062\,
            I => \dataRead3_14\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__20059\,
            I => \dataRead3_14\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__20056\,
            I => \dataRead3_14\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__20049\,
            I => \N__20044\
        );

    \I__3100\ : InMux
    port map (
            O => \N__20048\,
            I => \N__20041\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__20047\,
            I => \N__20038\
        );

    \I__3098\ : InMux
    port map (
            O => \N__20044\,
            I => \N__20035\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__20041\,
            I => \N__20032\
        );

    \I__3096\ : InMux
    port map (
            O => \N__20038\,
            I => \N__20029\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__20035\,
            I => \N__20024\
        );

    \I__3094\ : Span4Mux_h
    port map (
            O => \N__20032\,
            I => \N__20024\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__20029\,
            I => \dataRead2_14\
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__20024\,
            I => \dataRead2_14\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__20019\,
            I => \N__20016\
        );

    \I__3090\ : InMux
    port map (
            O => \N__20016\,
            I => \N__20013\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__20013\,
            I => \N__20009\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__20012\,
            I => \N__20005\
        );

    \I__3087\ : Span4Mux_v
    port map (
            O => \N__20009\,
            I => \N__20002\
        );

    \I__3086\ : InMux
    port map (
            O => \N__20008\,
            I => \N__19999\
        );

    \I__3085\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19996\
        );

    \I__3084\ : Span4Mux_h
    port map (
            O => \N__20002\,
            I => \N__19993\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__19999\,
            I => \dataRead5_13\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__19996\,
            I => \dataRead5_13\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__19993\,
            I => \dataRead5_13\
        );

    \I__3080\ : InMux
    port map (
            O => \N__19986\,
            I => \N__19983\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__19983\,
            I => \N__19980\
        );

    \I__3078\ : Span4Mux_v
    port map (
            O => \N__19980\,
            I => \N__19977\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__19977\,
            I => \QuadInstance2.Quad_RNO_0_2_13\
        );

    \I__3076\ : InMux
    port map (
            O => \N__19974\,
            I => \N__19970\
        );

    \I__3075\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19967\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__19970\,
            I => \N__19964\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__19967\,
            I => \N__19961\
        );

    \I__3072\ : Span4Mux_v
    port map (
            O => \N__19964\,
            I => \N__19957\
        );

    \I__3071\ : Span4Mux_h
    port map (
            O => \N__19961\,
            I => \N__19954\
        );

    \I__3070\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19951\
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__19957\,
            I => \dataRead2_13\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__19954\,
            I => \dataRead2_13\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__19951\,
            I => \dataRead2_13\
        );

    \I__3066\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19941\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__19941\,
            I => \QuadInstance3.Quad_RNO_0_3_13\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__3063\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19932\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__19932\,
            I => \N__19929\
        );

    \I__3061\ : Span4Mux_v
    port map (
            O => \N__19929\,
            I => \N__19925\
        );

    \I__3060\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19922\
        );

    \I__3059\ : Sp12to4
    port map (
            O => \N__19925\,
            I => \N__19918\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__19922\,
            I => \N__19915\
        );

    \I__3057\ : InMux
    port map (
            O => \N__19921\,
            I => \N__19912\
        );

    \I__3056\ : Odrv12
    port map (
            O => \N__19918\,
            I => \dataRead3_13\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__19915\,
            I => \dataRead3_13\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__19912\,
            I => \dataRead3_13\
        );

    \I__3053\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19902\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__19902\,
            I => \QuadInstance3.Quad_RNO_0_3_12\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__19899\,
            I => \N__19896\
        );

    \I__3050\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19893\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__19893\,
            I => \QuadInstance3.Quad_RNO_0_3_8\
        );

    \I__3048\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19887\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__19887\,
            I => \N__19884\
        );

    \I__3046\ : Span4Mux_h
    port map (
            O => \N__19884\,
            I => \N__19881\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__19881\,
            I => \QuadInstance7.Quad_RNO_0_7_7\
        );

    \I__3044\ : InMux
    port map (
            O => \N__19878\,
            I => \N__19875\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__19875\,
            I => \N__19872\
        );

    \I__3042\ : Odrv12
    port map (
            O => \N__19872\,
            I => \QuadInstance2.Quad_RNO_0_2_11\
        );

    \I__3041\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19866\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__19866\,
            I => \QuadInstance5.Quad_RNO_0_5_10\
        );

    \I__3039\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19860\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__19860\,
            I => \QuadInstance5.Quad_RNO_0_5_11\
        );

    \I__3037\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__19854\,
            I => \N__19851\
        );

    \I__3035\ : Span4Mux_h
    port map (
            O => \N__19851\,
            I => \N__19848\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__19848\,
            I => \QuadInstance2.Quad_RNO_0_2_8\
        );

    \I__3033\ : InMux
    port map (
            O => \N__19845\,
            I => \N__19842\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__19842\,
            I => \N__19839\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__19839\,
            I => \QuadInstance3.Quad_RNO_0_3_9\
        );

    \I__3030\ : InMux
    port map (
            O => \N__19836\,
            I => \N__19833\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__19833\,
            I => \N__19830\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__19827\,
            I => \QuadInstance7.Quad_RNO_0_7_9\
        );

    \I__3026\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__19821\,
            I => \N__19818\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__19818\,
            I => \QuadInstance5.Quad_RNO_0_5_8\
        );

    \I__3023\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__19812\,
            I => \N__19809\
        );

    \I__3021\ : Span4Mux_v
    port map (
            O => \N__19809\,
            I => \N__19806\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__19806\,
            I => \QuadInstance3.Quad_RNO_0_3_3\
        );

    \I__3019\ : InMux
    port map (
            O => \N__19803\,
            I => \N__19800\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__19800\,
            I => \N__19797\
        );

    \I__3017\ : Odrv12
    port map (
            O => \N__19797\,
            I => \QuadInstance2.Quad_RNO_0_2_7\
        );

    \I__3016\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19791\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__19788\,
            I => \QuadInstance3.Quad_RNO_0_3_7\
        );

    \I__3013\ : InMux
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__19782\,
            I => \QuadInstance5.Quad_RNO_0_5_7\
        );

    \I__3011\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19776\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__19776\,
            I => \N__19773\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__19773\,
            I => \QuadInstance3.Quad_RNO_0_3_5\
        );

    \I__3008\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__19767\,
            I => \N__19764\
        );

    \I__3006\ : Span4Mux_h
    port map (
            O => \N__19764\,
            I => \N__19761\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__19761\,
            I => \QuadInstance2.Quad_RNO_0_2_6\
        );

    \I__3004\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__19755\,
            I => \N__19752\
        );

    \I__3002\ : Span4Mux_h
    port map (
            O => \N__19752\,
            I => \N__19749\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__19749\,
            I => \QuadInstance7.Quad_RNO_0_7_2\
        );

    \I__3000\ : InMux
    port map (
            O => \N__19746\,
            I => \N__19743\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__19743\,
            I => \N__19740\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__19740\,
            I => \N__19737\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__19737\,
            I => \QuadInstance2.Quad_RNO_0_2_3\
        );

    \I__2996\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19731\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__19731\,
            I => \QuadInstance5.Quad_RNO_0_5_4\
        );

    \I__2994\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19725\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__19725\,
            I => \QuadInstance5.Quad_RNO_0_5_6\
        );

    \I__2992\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__19719\,
            I => \N__19716\
        );

    \I__2990\ : Span4Mux_h
    port map (
            O => \N__19716\,
            I => \N__19713\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__19713\,
            I => \QuadInstance7.Quad_RNO_0_7_6\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__19710\,
            I => \PWMInstance6.un1_periodCounter12_1_0_a2_0_0_cascade_\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__19707\,
            I => \PWMInstance6.un1_periodCounter12_1_0_a2_0_12_cascade_\
        );

    \I__2986\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19701\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__19701\,
            I => \PWMInstance6.un1_periodCounter12_1_0_a2_0_10\
        );

    \I__2984\ : InMux
    port map (
            O => \N__19698\,
            I => \N__19695\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__19695\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_2\
        );

    \I__2982\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19689\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__19689\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_3\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__19686\,
            I => \N__19683\
        );

    \I__2979\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19680\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__19680\,
            I => \PWMInstance6.PWMPulseWidthCountZ0Z_4\
        );

    \I__2977\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19674\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__19674\,
            I => \N__19671\
        );

    \I__2975\ : Span4Mux_v
    port map (
            O => \N__19671\,
            I => \N__19668\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__19668\,
            I => \QuadInstance2.Quad_RNO_0_2_2\
        );

    \I__2973\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19662\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__19662\,
            I => \N__19659\
        );

    \I__2971\ : Span4Mux_h
    port map (
            O => \N__19659\,
            I => \N__19656\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__19656\,
            I => \QuadInstance3.Quad_RNO_0_3_2\
        );

    \I__2969\ : CEMux
    port map (
            O => \N__19653\,
            I => \N__19646\
        );

    \I__2968\ : CEMux
    port map (
            O => \N__19652\,
            I => \N__19643\
        );

    \I__2967\ : CEMux
    port map (
            O => \N__19651\,
            I => \N__19640\
        );

    \I__2966\ : CEMux
    port map (
            O => \N__19650\,
            I => \N__19636\
        );

    \I__2965\ : CEMux
    port map (
            O => \N__19649\,
            I => \N__19632\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19627\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__19643\,
            I => \N__19627\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__19640\,
            I => \N__19624\
        );

    \I__2961\ : CEMux
    port map (
            O => \N__19639\,
            I => \N__19621\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__19636\,
            I => \N__19618\
        );

    \I__2959\ : CEMux
    port map (
            O => \N__19635\,
            I => \N__19615\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__19632\,
            I => \N__19612\
        );

    \I__2957\ : Span4Mux_v
    port map (
            O => \N__19627\,
            I => \N__19609\
        );

    \I__2956\ : Span4Mux_v
    port map (
            O => \N__19624\,
            I => \N__19606\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19603\
        );

    \I__2954\ : Span4Mux_h
    port map (
            O => \N__19618\,
            I => \N__19598\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__19615\,
            I => \N__19598\
        );

    \I__2952\ : Span4Mux_h
    port map (
            O => \N__19612\,
            I => \N__19594\
        );

    \I__2951\ : Span4Mux_h
    port map (
            O => \N__19609\,
            I => \N__19587\
        );

    \I__2950\ : Span4Mux_h
    port map (
            O => \N__19606\,
            I => \N__19587\
        );

    \I__2949\ : Span4Mux_v
    port map (
            O => \N__19603\,
            I => \N__19587\
        );

    \I__2948\ : Span4Mux_h
    port map (
            O => \N__19598\,
            I => \N__19584\
        );

    \I__2947\ : CEMux
    port map (
            O => \N__19597\,
            I => \N__19581\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__19594\,
            I => \PWMInstance5.pwmWrite_0_5\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__19587\,
            I => \PWMInstance5.pwmWrite_0_5\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__19584\,
            I => \PWMInstance5.pwmWrite_0_5\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__19581\,
            I => \PWMInstance5.pwmWrite_0_5\
        );

    \I__2942\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19562\
        );

    \I__2941\ : InMux
    port map (
            O => \N__19571\,
            I => \N__19562\
        );

    \I__2940\ : InMux
    port map (
            O => \N__19570\,
            I => \N__19562\
        );

    \I__2939\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19559\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__19562\,
            I => \PWMInstance5.clkCountZ0Z_1\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__19559\,
            I => \PWMInstance5.clkCountZ0Z_1\
        );

    \I__2936\ : InMux
    port map (
            O => \N__19554\,
            I => \N__19542\
        );

    \I__2935\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19542\
        );

    \I__2934\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19542\
        );

    \I__2933\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19542\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__19542\,
            I => \PWMInstance5.clkCountZ0Z_0\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__19539\,
            I => \N__19535\
        );

    \I__2930\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19532\
        );

    \I__2929\ : InMux
    port map (
            O => \N__19535\,
            I => \N__19529\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__19532\,
            I => \PWMInstance5.periodCounter12\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__19529\,
            I => \PWMInstance5.periodCounter12\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__19524\,
            I => \N__19520\
        );

    \I__2925\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19516\
        );

    \I__2924\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19513\
        );

    \I__2923\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19510\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__19516\,
            I => \PWMInstance5.periodCounterZ0Z_15\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__19513\,
            I => \PWMInstance5.periodCounterZ0Z_15\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__19510\,
            I => \PWMInstance5.periodCounterZ0Z_15\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__19503\,
            I => \N__19498\
        );

    \I__2918\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19495\
        );

    \I__2917\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19492\
        );

    \I__2916\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19489\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__19495\,
            I => \PWMInstance5.periodCounterZ0Z_1\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__19492\,
            I => \PWMInstance5.periodCounterZ0Z_1\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__19489\,
            I => \PWMInstance5.periodCounterZ0Z_1\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__19482\,
            I => \PWMInstance5.periodCounter12_cascade_\
        );

    \I__2911\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19476\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__19476\,
            I => \N__19473\
        );

    \I__2909\ : Odrv4
    port map (
            O => \N__19473\,
            I => \PWMInstance5.un1_periodCounter12_1_0_a2_0_9\
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__19470\,
            I => \PWMInstance5.un1_periodCounter12_1_0_a2_0_14_cascade_\
        );

    \I__2907\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__19464\,
            I => \PWMInstance5.un1_periodCounter12_1_0_a2_0_12\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__19461\,
            I => \N__19458\
        );

    \I__2904\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19455\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__19455\,
            I => \N__19447\
        );

    \I__2902\ : InMux
    port map (
            O => \N__19454\,
            I => \N__19442\
        );

    \I__2901\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19442\
        );

    \I__2900\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19439\
        );

    \I__2899\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19436\
        );

    \I__2898\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19433\
        );

    \I__2897\ : Span12Mux_v
    port map (
            O => \N__19447\,
            I => \N__19430\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__19442\,
            I => \PWMInstance5.out_0_sqmuxa\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__19439\,
            I => \PWMInstance5.out_0_sqmuxa\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__19436\,
            I => \PWMInstance5.out_0_sqmuxa\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__19433\,
            I => \PWMInstance5.out_0_sqmuxa\
        );

    \I__2892\ : Odrv12
    port map (
            O => \N__19430\,
            I => \PWMInstance5.out_0_sqmuxa\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__19419\,
            I => \N__19416\
        );

    \I__2890\ : InMux
    port map (
            O => \N__19416\,
            I => \N__19411\
        );

    \I__2889\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19408\
        );

    \I__2888\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19405\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__19411\,
            I => \N__19402\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__19408\,
            I => \PWMInstance5.periodCounterZ0Z_9\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__19405\,
            I => \PWMInstance5.periodCounterZ0Z_9\
        );

    \I__2884\ : Odrv12
    port map (
            O => \N__19402\,
            I => \PWMInstance5.periodCounterZ0Z_9\
        );

    \I__2883\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19390\
        );

    \I__2882\ : CascadeMux
    port map (
            O => \N__19394\,
            I => \N__19387\
        );

    \I__2881\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19384\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__19390\,
            I => \N__19381\
        );

    \I__2879\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19378\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__19384\,
            I => \PWMInstance5.periodCounterZ0Z_5\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__19381\,
            I => \PWMInstance5.periodCounterZ0Z_5\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__19378\,
            I => \PWMInstance5.periodCounterZ0Z_5\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__19371\,
            I => \N__19366\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__19370\,
            I => \N__19363\
        );

    \I__2873\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19360\
        );

    \I__2872\ : InMux
    port map (
            O => \N__19366\,
            I => \N__19357\
        );

    \I__2871\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19354\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__19360\,
            I => \PWMInstance5.periodCounterZ0Z_11\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__19357\,
            I => \PWMInstance5.periodCounterZ0Z_11\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__19354\,
            I => \PWMInstance5.periodCounterZ0Z_11\
        );

    \I__2867\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19342\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__19346\,
            I => \N__19339\
        );

    \I__2865\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19336\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__19342\,
            I => \N__19333\
        );

    \I__2863\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19330\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__19336\,
            I => \PWMInstance5.periodCounterZ0Z_3\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__19333\,
            I => \PWMInstance5.periodCounterZ0Z_3\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__19330\,
            I => \PWMInstance5.periodCounterZ0Z_3\
        );

    \I__2859\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19320\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__19320\,
            I => \PWMInstance5.un1_periodCounter12_1_0_a2_0_10\
        );

    \I__2857\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19312\
        );

    \I__2856\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19309\
        );

    \I__2855\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19306\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__19312\,
            I => \PWMInstance5.periodCounterZ0Z_16\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__19309\,
            I => \PWMInstance5.periodCounterZ0Z_16\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__19306\,
            I => \PWMInstance5.periodCounterZ0Z_16\
        );

    \I__2851\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19294\
        );

    \I__2850\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19291\
        );

    \I__2849\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19288\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__19294\,
            I => \N__19285\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__19291\,
            I => \PWMInstance5.periodCounterZ0Z_7\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__19288\,
            I => \PWMInstance5.periodCounterZ0Z_7\
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__19285\,
            I => \PWMInstance5.periodCounterZ0Z_7\
        );

    \I__2844\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19275\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__19275\,
            I => \PWMInstance5.un1_periodCounter12_1_0_a2_0_6\
        );

    \I__2842\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19269\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__19269\,
            I => \N__19266\
        );

    \I__2840\ : Span4Mux_h
    port map (
            O => \N__19266\,
            I => \N__19263\
        );

    \I__2839\ : Span4Mux_v
    port map (
            O => \N__19263\,
            I => \N__19260\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__19260\,
            I => \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_4\
        );

    \I__2837\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19252\
        );

    \I__2836\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19249\
        );

    \I__2835\ : InMux
    port map (
            O => \N__19255\,
            I => \N__19246\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__19252\,
            I => \PWMInstance5.periodCounterZ0Z_2\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__19249\,
            I => \PWMInstance5.periodCounterZ0Z_2\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__19246\,
            I => \PWMInstance5.periodCounterZ0Z_2\
        );

    \I__2831\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19234\
        );

    \I__2830\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19231\
        );

    \I__2829\ : InMux
    port map (
            O => \N__19237\,
            I => \N__19228\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__19234\,
            I => \PWMInstance5.periodCounterZ0Z_14\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__19231\,
            I => \PWMInstance5.periodCounterZ0Z_14\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__19228\,
            I => \PWMInstance5.periodCounterZ0Z_14\
        );

    \I__2825\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19216\
        );

    \I__2824\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19213\
        );

    \I__2823\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19210\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__19216\,
            I => \PWMInstance5.periodCounterZ0Z_12\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__19213\,
            I => \PWMInstance5.periodCounterZ0Z_12\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__19210\,
            I => \PWMInstance5.periodCounterZ0Z_12\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__19203\,
            I => \PWMInstance5.un1_periodCounter12_1_0_a2_0_0_cascade_\
        );

    \I__2818\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19195\
        );

    \I__2817\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19190\
        );

    \I__2816\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19190\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__19195\,
            I => \PWMInstance5.periodCounterZ0Z_4\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__19190\,
            I => \PWMInstance5.periodCounterZ0Z_4\
        );

    \I__2813\ : InMux
    port map (
            O => \N__19185\,
            I => \N__19182\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__19182\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_4\
        );

    \I__2811\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19176\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__19176\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_5\
        );

    \I__2809\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19168\
        );

    \I__2808\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19163\
        );

    \I__2807\ : InMux
    port map (
            O => \N__19171\,
            I => \N__19163\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__19168\,
            I => \PWMInstance5.periodCounterZ0Z_10\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__19163\,
            I => \PWMInstance5.periodCounterZ0Z_10\
        );

    \I__2804\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19155\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__19155\,
            I => \N__19152\
        );

    \I__2802\ : Span4Mux_h
    port map (
            O => \N__19152\,
            I => \N__19149\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__19149\,
            I => \N__19146\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__19146\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_10\
        );

    \I__2799\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__19140\,
            I => \N__19137\
        );

    \I__2797\ : Span4Mux_h
    port map (
            O => \N__19137\,
            I => \N__19134\
        );

    \I__2796\ : Span4Mux_v
    port map (
            O => \N__19134\,
            I => \N__19131\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__19131\,
            I => \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_4\
        );

    \I__2794\ : InMux
    port map (
            O => \N__19128\,
            I => \N__19125\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__19125\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_11\
        );

    \I__2792\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19119\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__19119\,
            I => \N__19116\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__19116\,
            I => \N__19113\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__19113\,
            I => \N__19110\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__19110\,
            I => \PWMInstance5.un1_periodCounter12_1_0_a2_0\
        );

    \I__2787\ : InMux
    port map (
            O => \N__19107\,
            I => \N__19104\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__19104\,
            I => \N__19101\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__19101\,
            I => \QuadInstance3.Quad_RNIBRAL1Z0Z_4\
        );

    \I__2784\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19095\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__19095\,
            I => \N__19092\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__19092\,
            I => \QuadInstance3.Quad_RNIS50J1Z0Z_14\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__19089\,
            I => \N__19085\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__19088\,
            I => \N__19082\
        );

    \I__2779\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19077\
        );

    \I__2778\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19077\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__19077\,
            I => \QuadInstance3.delayedCh_BZ0Z_2\
        );

    \I__2776\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19071\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__19071\,
            I => \QuadInstance3.delayedCh_AZ0Z_2\
        );

    \I__2774\ : InMux
    port map (
            O => \N__19068\,
            I => \N__19063\
        );

    \I__2773\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19058\
        );

    \I__2772\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19058\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__19063\,
            I => \QuadInstance3.delayedCh_AZ0Z_1\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__19058\,
            I => \QuadInstance3.delayedCh_AZ0Z_1\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__19053\,
            I => \N__19050\
        );

    \I__2768\ : InMux
    port map (
            O => \N__19050\,
            I => \N__19047\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__19047\,
            I => \N__19044\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__19044\,
            I => \QuadInstance3.Quad_RNIEUAL1Z0Z_7\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__19041\,
            I => \N__19036\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__19040\,
            I => \N__19031\
        );

    \I__2763\ : InMux
    port map (
            O => \N__19039\,
            I => \N__19015\
        );

    \I__2762\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19015\
        );

    \I__2761\ : InMux
    port map (
            O => \N__19035\,
            I => \N__19015\
        );

    \I__2760\ : InMux
    port map (
            O => \N__19034\,
            I => \N__19008\
        );

    \I__2759\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19008\
        );

    \I__2758\ : InMux
    port map (
            O => \N__19030\,
            I => \N__19008\
        );

    \I__2757\ : InMux
    port map (
            O => \N__19029\,
            I => \N__19001\
        );

    \I__2756\ : InMux
    port map (
            O => \N__19028\,
            I => \N__19001\
        );

    \I__2755\ : InMux
    port map (
            O => \N__19027\,
            I => \N__19001\
        );

    \I__2754\ : InMux
    port map (
            O => \N__19026\,
            I => \N__18994\
        );

    \I__2753\ : InMux
    port map (
            O => \N__19025\,
            I => \N__18994\
        );

    \I__2752\ : InMux
    port map (
            O => \N__19024\,
            I => \N__18994\
        );

    \I__2751\ : InMux
    port map (
            O => \N__19023\,
            I => \N__18989\
        );

    \I__2750\ : InMux
    port map (
            O => \N__19022\,
            I => \N__18989\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__19015\,
            I => \QuadInstance3.un1_count_enable_i_a2_0_1\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__19008\,
            I => \QuadInstance3.un1_count_enable_i_a2_0_1\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__19001\,
            I => \QuadInstance3.un1_count_enable_i_a2_0_1\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__18994\,
            I => \QuadInstance3.un1_count_enable_i_a2_0_1\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__18989\,
            I => \QuadInstance3.un1_count_enable_i_a2_0_1\
        );

    \I__2744\ : InMux
    port map (
            O => \N__18978\,
            I => \N__18968\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__18977\,
            I => \N__18965\
        );

    \I__2742\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18961\
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__18975\,
            I => \N__18958\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__18974\,
            I => \N__18955\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__18973\,
            I => \N__18951\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__18972\,
            I => \N__18942\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__18971\,
            I => \N__18939\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__18968\,
            I => \N__18936\
        );

    \I__2735\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18931\
        );

    \I__2734\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18931\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18928\
        );

    \I__2732\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18925\
        );

    \I__2731\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18914\
        );

    \I__2730\ : InMux
    port map (
            O => \N__18954\,
            I => \N__18914\
        );

    \I__2729\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18914\
        );

    \I__2728\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18914\
        );

    \I__2727\ : InMux
    port map (
            O => \N__18949\,
            I => \N__18914\
        );

    \I__2726\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18901\
        );

    \I__2725\ : InMux
    port map (
            O => \N__18947\,
            I => \N__18901\
        );

    \I__2724\ : InMux
    port map (
            O => \N__18946\,
            I => \N__18901\
        );

    \I__2723\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18901\
        );

    \I__2722\ : InMux
    port map (
            O => \N__18942\,
            I => \N__18901\
        );

    \I__2721\ : InMux
    port map (
            O => \N__18939\,
            I => \N__18901\
        );

    \I__2720\ : Odrv12
    port map (
            O => \N__18936\,
            I => \QuadInstance3.count_enable\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__18931\,
            I => \QuadInstance3.count_enable\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__18928\,
            I => \QuadInstance3.count_enable\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__18925\,
            I => \QuadInstance3.count_enable\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__18914\,
            I => \QuadInstance3.count_enable\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__18901\,
            I => \QuadInstance3.count_enable\
        );

    \I__2714\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18885\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__18885\,
            I => \N__18882\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__18882\,
            I => \QuadInstance3.un1_Quad_axb_15\
        );

    \I__2711\ : InMux
    port map (
            O => \N__18879\,
            I => \N__18876\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__18876\,
            I => \N__18873\
        );

    \I__2709\ : Span4Mux_v
    port map (
            O => \N__18873\,
            I => \N__18870\
        );

    \I__2708\ : Span4Mux_v
    port map (
            O => \N__18870\,
            I => \N__18867\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__18867\,
            I => \QuadInstance3.delayedCh_BZ0Z_0\
        );

    \I__2706\ : InMux
    port map (
            O => \N__18864\,
            I => \N__18860\
        );

    \I__2705\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18857\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__18860\,
            I => \QuadInstance3.delayedCh_BZ0Z_1\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__18857\,
            I => \QuadInstance3.delayedCh_BZ0Z_1\
        );

    \I__2702\ : InMux
    port map (
            O => \N__18852\,
            I => \QuadInstance3.un1_Quad_cry_13\
        );

    \I__2701\ : InMux
    port map (
            O => \N__18849\,
            I => \QuadInstance3.un1_Quad_cry_14\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__18846\,
            I => \QuadInstance3.count_enable_cascade_\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__18843\,
            I => \N__18840\
        );

    \I__2698\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18837\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__18837\,
            I => \N__18834\
        );

    \I__2696\ : Odrv4
    port map (
            O => \N__18834\,
            I => \QuadInstance3.Quad_RNI8OAL1Z0Z_1\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__18831\,
            I => \QuadInstance3.un1_count_enable_i_a2_0_1_cascade_\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__18828\,
            I => \N__18825\
        );

    \I__2693\ : InMux
    port map (
            O => \N__18825\,
            I => \N__18822\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__18822\,
            I => \N__18819\
        );

    \I__2691\ : Odrv4
    port map (
            O => \N__18819\,
            I => \QuadInstance3.Quad_RNI9PAL1Z0Z_2\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__18816\,
            I => \N__18813\
        );

    \I__2689\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18810\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__18810\,
            I => \QuadInstance3.Quad_RNIO10J1Z0Z_10\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__18807\,
            I => \N__18804\
        );

    \I__2686\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18801\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__18801\,
            I => \QuadInstance3.Quad_RNIFVAL1Z0Z_8\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__18798\,
            I => \N__18795\
        );

    \I__2683\ : InMux
    port map (
            O => \N__18795\,
            I => \N__18792\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__18792\,
            I => \QuadInstance3.Quad_RNIG0BL1Z0Z_9\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__18789\,
            I => \N__18786\
        );

    \I__2680\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18783\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__18783\,
            I => \N__18780\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__18780\,
            I => \QuadInstance3.Quad_RNICSAL1Z0Z_5\
        );

    \I__2677\ : InMux
    port map (
            O => \N__18777\,
            I => \QuadInstance3.un1_Quad_cry_4\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__18774\,
            I => \N__18771\
        );

    \I__2675\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18768\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__18768\,
            I => \N__18765\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__18765\,
            I => \QuadInstance3.Quad_RNIDTAL1Z0Z_6\
        );

    \I__2672\ : InMux
    port map (
            O => \N__18762\,
            I => \QuadInstance3.un1_Quad_cry_5\
        );

    \I__2671\ : InMux
    port map (
            O => \N__18759\,
            I => \QuadInstance3.un1_Quad_cry_6\
        );

    \I__2670\ : InMux
    port map (
            O => \N__18756\,
            I => \bfn_10_9_0_\
        );

    \I__2669\ : InMux
    port map (
            O => \N__18753\,
            I => \QuadInstance3.un1_Quad_cry_8\
        );

    \I__2668\ : InMux
    port map (
            O => \N__18750\,
            I => \QuadInstance3.un1_Quad_cry_9\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__18747\,
            I => \N__18744\
        );

    \I__2666\ : InMux
    port map (
            O => \N__18744\,
            I => \N__18741\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__18741\,
            I => \QuadInstance3.Quad_RNIP20J1Z0Z_11\
        );

    \I__2664\ : InMux
    port map (
            O => \N__18738\,
            I => \QuadInstance3.un1_Quad_cry_10\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__18735\,
            I => \N__18732\
        );

    \I__2662\ : InMux
    port map (
            O => \N__18732\,
            I => \N__18729\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__18729\,
            I => \QuadInstance3.Quad_RNIQ30J1Z0Z_12\
        );

    \I__2660\ : InMux
    port map (
            O => \N__18726\,
            I => \QuadInstance3.un1_Quad_cry_11\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__18723\,
            I => \N__18720\
        );

    \I__2658\ : InMux
    port map (
            O => \N__18720\,
            I => \N__18717\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__18717\,
            I => \QuadInstance3.Quad_RNIR40J1Z0Z_13\
        );

    \I__2656\ : InMux
    port map (
            O => \N__18714\,
            I => \QuadInstance3.un1_Quad_cry_12\
        );

    \I__2655\ : InMux
    port map (
            O => \N__18711\,
            I => \N__18708\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__18708\,
            I => \QuadInstance5.Quad_RNIBDQ82Z0Z_13\
        );

    \I__2653\ : InMux
    port map (
            O => \N__18705\,
            I => \N__18702\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__18702\,
            I => \QuadInstance5.Quad_RNO_0_5_13\
        );

    \I__2651\ : InMux
    port map (
            O => \N__18699\,
            I => \QuadInstance5.un1_Quad_cry_12\
        );

    \I__2650\ : InMux
    port map (
            O => \N__18696\,
            I => \N__18693\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__18693\,
            I => \QuadInstance5.Quad_RNICEQ82Z0Z_14\
        );

    \I__2648\ : InMux
    port map (
            O => \N__18690\,
            I => \N__18687\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__18687\,
            I => \QuadInstance5.Quad_RNO_0_5_14\
        );

    \I__2646\ : InMux
    port map (
            O => \N__18684\,
            I => \QuadInstance5.un1_Quad_cry_13\
        );

    \I__2645\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18678\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__18678\,
            I => \QuadInstance5.un1_Quad_axb_15\
        );

    \I__2643\ : InMux
    port map (
            O => \N__18675\,
            I => \QuadInstance5.un1_Quad_cry_14\
        );

    \I__2642\ : InMux
    port map (
            O => \N__18672\,
            I => \QuadInstance3.un1_Quad_cry_0\
        );

    \I__2641\ : InMux
    port map (
            O => \N__18669\,
            I => \QuadInstance3.un1_Quad_cry_1\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__18666\,
            I => \N__18663\
        );

    \I__2639\ : InMux
    port map (
            O => \N__18663\,
            I => \N__18660\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__18660\,
            I => \N__18657\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__18657\,
            I => \QuadInstance3.Quad_RNIAQAL1Z0Z_3\
        );

    \I__2636\ : InMux
    port map (
            O => \N__18654\,
            I => \QuadInstance3.un1_Quad_cry_2\
        );

    \I__2635\ : InMux
    port map (
            O => \N__18651\,
            I => \QuadInstance3.un1_Quad_cry_3\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__18648\,
            I => \N__18645\
        );

    \I__2633\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18642\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__18642\,
            I => \QuadInstance5.Quad_RNIR1LI2Z0Z_4\
        );

    \I__2631\ : InMux
    port map (
            O => \N__18639\,
            I => \QuadInstance5.un1_Quad_cry_3\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__18636\,
            I => \N__18633\
        );

    \I__2629\ : InMux
    port map (
            O => \N__18633\,
            I => \N__18630\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__18630\,
            I => \QuadInstance5.Quad_RNIS2LI2Z0Z_5\
        );

    \I__2627\ : InMux
    port map (
            O => \N__18627\,
            I => \QuadInstance5.un1_Quad_cry_4\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__18624\,
            I => \N__18621\
        );

    \I__2625\ : InMux
    port map (
            O => \N__18621\,
            I => \N__18618\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__18618\,
            I => \QuadInstance5.Quad_RNIT3LI2Z0Z_6\
        );

    \I__2623\ : InMux
    port map (
            O => \N__18615\,
            I => \QuadInstance5.un1_Quad_cry_5\
        );

    \I__2622\ : InMux
    port map (
            O => \N__18612\,
            I => \N__18609\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__18609\,
            I => \QuadInstance5.Quad_RNIU4LI2Z0Z_7\
        );

    \I__2620\ : InMux
    port map (
            O => \N__18606\,
            I => \QuadInstance5.un1_Quad_cry_6\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__18603\,
            I => \N__18600\
        );

    \I__2618\ : InMux
    port map (
            O => \N__18600\,
            I => \N__18597\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__18597\,
            I => \QuadInstance5.Quad_RNIV5LI2Z0Z_8\
        );

    \I__2616\ : InMux
    port map (
            O => \N__18594\,
            I => \bfn_10_7_0_\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__18591\,
            I => \N__18588\
        );

    \I__2614\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18585\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__18585\,
            I => \N__18582\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__18582\,
            I => \QuadInstance5.Quad_RNI07LI2Z0Z_9\
        );

    \I__2611\ : InMux
    port map (
            O => \N__18579\,
            I => \QuadInstance5.un1_Quad_cry_8\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__18576\,
            I => \N__18573\
        );

    \I__2609\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18570\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__18570\,
            I => \QuadInstance5.Quad_RNI8AQ82Z0Z_10\
        );

    \I__2607\ : InMux
    port map (
            O => \N__18567\,
            I => \QuadInstance5.un1_Quad_cry_9\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__18564\,
            I => \N__18561\
        );

    \I__2605\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18558\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__18558\,
            I => \QuadInstance5.Quad_RNI9BQ82Z0Z_11\
        );

    \I__2603\ : InMux
    port map (
            O => \N__18555\,
            I => \QuadInstance5.un1_Quad_cry_10\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__18552\,
            I => \N__18549\
        );

    \I__2601\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18546\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__18546\,
            I => \QuadInstance5.Quad_RNIACQ82Z0Z_12\
        );

    \I__2599\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18540\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__18540\,
            I => \QuadInstance5.Quad_RNO_0_5_12\
        );

    \I__2597\ : InMux
    port map (
            O => \N__18537\,
            I => \QuadInstance5.un1_Quad_cry_11\
        );

    \I__2596\ : InMux
    port map (
            O => \N__18534\,
            I => \N__18531\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__18531\,
            I => \N__18526\
        );

    \I__2594\ : InMux
    port map (
            O => \N__18530\,
            I => \N__18523\
        );

    \I__2593\ : InMux
    port map (
            O => \N__18529\,
            I => \N__18520\
        );

    \I__2592\ : Span4Mux_v
    port map (
            O => \N__18526\,
            I => \N__18508\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__18523\,
            I => \N__18508\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__18520\,
            I => \N__18508\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__18519\,
            I => \N__18500\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__18518\,
            I => \N__18496\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__18517\,
            I => \N__18493\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__18516\,
            I => \N__18488\
        );

    \I__2585\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18485\
        );

    \I__2584\ : Span4Mux_h
    port map (
            O => \N__18508\,
            I => \N__18482\
        );

    \I__2583\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18473\
        );

    \I__2582\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18473\
        );

    \I__2581\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18473\
        );

    \I__2580\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18473\
        );

    \I__2579\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18456\
        );

    \I__2578\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18456\
        );

    \I__2577\ : InMux
    port map (
            O => \N__18499\,
            I => \N__18456\
        );

    \I__2576\ : InMux
    port map (
            O => \N__18496\,
            I => \N__18456\
        );

    \I__2575\ : InMux
    port map (
            O => \N__18493\,
            I => \N__18456\
        );

    \I__2574\ : InMux
    port map (
            O => \N__18492\,
            I => \N__18456\
        );

    \I__2573\ : InMux
    port map (
            O => \N__18491\,
            I => \N__18456\
        );

    \I__2572\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18456\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__18485\,
            I => \QuadInstance2.count_enable\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__18482\,
            I => \QuadInstance2.count_enable\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__18473\,
            I => \QuadInstance2.count_enable\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__18456\,
            I => \QuadInstance2.count_enable\
        );

    \I__2567\ : InMux
    port map (
            O => \N__18447\,
            I => \N__18443\
        );

    \I__2566\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18440\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__18443\,
            I => \QuadInstance5.delayedCh_BZ0Z_1\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__18440\,
            I => \QuadInstance5.delayedCh_BZ0Z_1\
        );

    \I__2563\ : InMux
    port map (
            O => \N__18435\,
            I => \N__18430\
        );

    \I__2562\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18427\
        );

    \I__2561\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18424\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__18430\,
            I => \QuadInstance5.delayedCh_AZ0Z_1\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__18427\,
            I => \QuadInstance5.delayedCh_AZ0Z_1\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__18424\,
            I => \QuadInstance5.delayedCh_AZ0Z_1\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__18417\,
            I => \N__18414\
        );

    \I__2556\ : InMux
    port map (
            O => \N__18414\,
            I => \N__18411\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__18411\,
            I => \QuadInstance5.delayedCh_AZ0Z_2\
        );

    \I__2554\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18404\
        );

    \I__2553\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18401\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__18404\,
            I => \QuadInstance5.delayedCh_BZ0Z_2\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__18401\,
            I => \QuadInstance5.delayedCh_BZ0Z_2\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__18396\,
            I => \QuadInstance5.count_enable_cascade_\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__18393\,
            I => \N__18389\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__18392\,
            I => \N__18384\
        );

    \I__2547\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18370\
        );

    \I__2546\ : InMux
    port map (
            O => \N__18388\,
            I => \N__18370\
        );

    \I__2545\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18370\
        );

    \I__2544\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18370\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__18383\,
            I => \N__18365\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__18382\,
            I => \N__18361\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__18381\,
            I => \N__18355\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__18380\,
            I => \N__18352\
        );

    \I__2539\ : CascadeMux
    port map (
            O => \N__18379\,
            I => \N__18348\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__18370\,
            I => \N__18345\
        );

    \I__2537\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18342\
        );

    \I__2536\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18331\
        );

    \I__2535\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18331\
        );

    \I__2534\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18331\
        );

    \I__2533\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18331\
        );

    \I__2532\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18331\
        );

    \I__2531\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18318\
        );

    \I__2530\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18318\
        );

    \I__2529\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18318\
        );

    \I__2528\ : InMux
    port map (
            O => \N__18352\,
            I => \N__18318\
        );

    \I__2527\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18318\
        );

    \I__2526\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18318\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__18345\,
            I => \QuadInstance5.count_enable\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__18342\,
            I => \QuadInstance5.count_enable\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__18331\,
            I => \QuadInstance5.count_enable\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__18318\,
            I => \QuadInstance5.count_enable\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__18309\,
            I => \N__18306\
        );

    \I__2520\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18303\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__18303\,
            I => \QuadInstance5.Quad_RNIOUKI2Z0Z_1\
        );

    \I__2518\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18297\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__18297\,
            I => \QuadInstance5.Quad_RNO_0_4_1\
        );

    \I__2516\ : InMux
    port map (
            O => \N__18294\,
            I => \QuadInstance5.un1_Quad_cry_0\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__18291\,
            I => \N__18288\
        );

    \I__2514\ : InMux
    port map (
            O => \N__18288\,
            I => \N__18285\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__18285\,
            I => \QuadInstance5.Quad_RNIPVKI2Z0Z_2\
        );

    \I__2512\ : InMux
    port map (
            O => \N__18282\,
            I => \QuadInstance5.un1_Quad_cry_1\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__18279\,
            I => \N__18276\
        );

    \I__2510\ : InMux
    port map (
            O => \N__18276\,
            I => \N__18273\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__18273\,
            I => \QuadInstance5.Quad_RNIQ0LI2Z0Z_3\
        );

    \I__2508\ : InMux
    port map (
            O => \N__18270\,
            I => \QuadInstance5.un1_Quad_cry_2\
        );

    \I__2507\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18264\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__18264\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_1\
        );

    \I__2505\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18258\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__18258\,
            I => \N__18255\
        );

    \I__2503\ : Span4Mux_h
    port map (
            O => \N__18255\,
            I => \N__18252\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__18252\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_7\
        );

    \I__2501\ : CEMux
    port map (
            O => \N__18249\,
            I => \N__18245\
        );

    \I__2500\ : CEMux
    port map (
            O => \N__18248\,
            I => \N__18242\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__18245\,
            I => \N__18239\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__18242\,
            I => \N__18236\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__18239\,
            I => \N__18228\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__18236\,
            I => \N__18228\
        );

    \I__2495\ : CEMux
    port map (
            O => \N__18235\,
            I => \N__18225\
        );

    \I__2494\ : CEMux
    port map (
            O => \N__18234\,
            I => \N__18222\
        );

    \I__2493\ : CEMux
    port map (
            O => \N__18233\,
            I => \N__18219\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__18228\,
            I => \PWMInstance0.pwmWrite_0_0\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__18225\,
            I => \PWMInstance0.pwmWrite_0_0\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__18222\,
            I => \PWMInstance0.pwmWrite_0_0\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__18219\,
            I => \PWMInstance0.pwmWrite_0_0\
        );

    \I__2488\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18207\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__18207\,
            I => \N__18204\
        );

    \I__2486\ : Odrv4
    port map (
            O => \N__18204\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_13\
        );

    \I__2485\ : InMux
    port map (
            O => \N__18201\,
            I => \N__18198\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__18198\,
            I => \N__18195\
        );

    \I__2483\ : Span12Mux_h
    port map (
            O => \N__18195\,
            I => \N__18192\
        );

    \I__2482\ : Odrv12
    port map (
            O => \N__18192\,
            I => \ch5_B_c\
        );

    \I__2481\ : InMux
    port map (
            O => \N__18189\,
            I => \N__18186\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__18186\,
            I => \N__18183\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__18183\,
            I => \QuadInstance5.delayedCh_BZ0Z_0\
        );

    \I__2478\ : InMux
    port map (
            O => \N__18180\,
            I => \PWMInstance5.un1_periodCounter_2_cry_11\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__18177\,
            I => \N__18174\
        );

    \I__2476\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18169\
        );

    \I__2475\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18166\
        );

    \I__2474\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18163\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__18169\,
            I => \N__18158\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__18166\,
            I => \N__18158\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__18163\,
            I => \PWMInstance5.periodCounterZ0Z_13\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__18158\,
            I => \PWMInstance5.periodCounterZ0Z_13\
        );

    \I__2469\ : InMux
    port map (
            O => \N__18153\,
            I => \PWMInstance5.un1_periodCounter_2_cry_12\
        );

    \I__2468\ : InMux
    port map (
            O => \N__18150\,
            I => \PWMInstance5.un1_periodCounter_2_cry_13\
        );

    \I__2467\ : InMux
    port map (
            O => \N__18147\,
            I => \PWMInstance5.un1_periodCounter_2_cry_14\
        );

    \I__2466\ : InMux
    port map (
            O => \N__18144\,
            I => \bfn_9_14_0_\
        );

    \I__2465\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18137\
        );

    \I__2464\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18134\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__18137\,
            I => \N__18130\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__18134\,
            I => \N__18127\
        );

    \I__2461\ : InMux
    port map (
            O => \N__18133\,
            I => \N__18124\
        );

    \I__2460\ : Span4Mux_h
    port map (
            O => \N__18130\,
            I => \N__18121\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__18127\,
            I => \N__18118\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__18124\,
            I => \PWMInstance0.periodCounterZ0Z_8\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__18121\,
            I => \PWMInstance0.periodCounterZ0Z_8\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__18118\,
            I => \PWMInstance0.periodCounterZ0Z_8\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__18111\,
            I => \N__18107\
        );

    \I__2454\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18104\
        );

    \I__2453\ : InMux
    port map (
            O => \N__18107\,
            I => \N__18101\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__18104\,
            I => \N__18097\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__18101\,
            I => \N__18094\
        );

    \I__2450\ : InMux
    port map (
            O => \N__18100\,
            I => \N__18091\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__18097\,
            I => \N__18088\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__18094\,
            I => \N__18085\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__18091\,
            I => \PWMInstance0.periodCounterZ0Z_6\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__18088\,
            I => \PWMInstance0.periodCounterZ0Z_6\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__18085\,
            I => \PWMInstance0.periodCounterZ0Z_6\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__18078\,
            I => \N__18074\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__18077\,
            I => \N__18071\
        );

    \I__2442\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18068\
        );

    \I__2441\ : InMux
    port map (
            O => \N__18071\,
            I => \N__18064\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__18068\,
            I => \N__18061\
        );

    \I__2439\ : InMux
    port map (
            O => \N__18067\,
            I => \N__18058\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__18064\,
            I => \N__18055\
        );

    \I__2437\ : Span4Mux_h
    port map (
            O => \N__18061\,
            I => \N__18052\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__18058\,
            I => \PWMInstance0.periodCounterZ0Z_13\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__18055\,
            I => \PWMInstance0.periodCounterZ0Z_13\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__18052\,
            I => \PWMInstance0.periodCounterZ0Z_13\
        );

    \I__2433\ : InMux
    port map (
            O => \N__18045\,
            I => \N__18042\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__18042\,
            I => \N__18039\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__18039\,
            I => \PWMInstance0.un1_periodCounter12_1_0_a2_0_9\
        );

    \I__2430\ : InMux
    port map (
            O => \N__18036\,
            I => \N__18029\
        );

    \I__2429\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18029\
        );

    \I__2428\ : InMux
    port map (
            O => \N__18034\,
            I => \N__18026\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__18029\,
            I => \N__18023\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__18026\,
            I => \N__18018\
        );

    \I__2425\ : Span4Mux_v
    port map (
            O => \N__18023\,
            I => \N__18018\
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__18018\,
            I => \PWMInstance0.periodCounterZ0Z_0\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__18015\,
            I => \N__18012\
        );

    \I__2422\ : InMux
    port map (
            O => \N__18012\,
            I => \N__18008\
        );

    \I__2421\ : InMux
    port map (
            O => \N__18011\,
            I => \N__18004\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__18008\,
            I => \N__18001\
        );

    \I__2419\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17998\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__18004\,
            I => \N__17993\
        );

    \I__2417\ : Span4Mux_v
    port map (
            O => \N__18001\,
            I => \N__17993\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__17998\,
            I => \PWMInstance0.periodCounterZ0Z_1\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__17993\,
            I => \PWMInstance0.periodCounterZ0Z_1\
        );

    \I__2414\ : InMux
    port map (
            O => \N__17988\,
            I => \N__17985\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__17985\,
            I => \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNOZ0\
        );

    \I__2412\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17979\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__17979\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_0\
        );

    \I__2410\ : InMux
    port map (
            O => \N__17976\,
            I => \PWMInstance5.un1_periodCounter_2_cry_2\
        );

    \I__2409\ : InMux
    port map (
            O => \N__17973\,
            I => \PWMInstance5.un1_periodCounter_2_cry_3\
        );

    \I__2408\ : InMux
    port map (
            O => \N__17970\,
            I => \PWMInstance5.un1_periodCounter_2_cry_4\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__17967\,
            I => \N__17963\
        );

    \I__2406\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17959\
        );

    \I__2405\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17954\
        );

    \I__2404\ : InMux
    port map (
            O => \N__17962\,
            I => \N__17954\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__17959\,
            I => \PWMInstance5.periodCounterZ0Z_6\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__17954\,
            I => \PWMInstance5.periodCounterZ0Z_6\
        );

    \I__2401\ : InMux
    port map (
            O => \N__17949\,
            I => \PWMInstance5.un1_periodCounter_2_cry_5\
        );

    \I__2400\ : InMux
    port map (
            O => \N__17946\,
            I => \PWMInstance5.un1_periodCounter_2_cry_6\
        );

    \I__2399\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17938\
        );

    \I__2398\ : InMux
    port map (
            O => \N__17942\,
            I => \N__17935\
        );

    \I__2397\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17932\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__17938\,
            I => \N__17929\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__17935\,
            I => \N__17926\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__17932\,
            I => \PWMInstance5.periodCounterZ0Z_8\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__17929\,
            I => \PWMInstance5.periodCounterZ0Z_8\
        );

    \I__2392\ : Odrv12
    port map (
            O => \N__17926\,
            I => \PWMInstance5.periodCounterZ0Z_8\
        );

    \I__2391\ : InMux
    port map (
            O => \N__17919\,
            I => \bfn_9_13_0_\
        );

    \I__2390\ : InMux
    port map (
            O => \N__17916\,
            I => \PWMInstance5.un1_periodCounter_2_cry_8\
        );

    \I__2389\ : InMux
    port map (
            O => \N__17913\,
            I => \PWMInstance5.un1_periodCounter_2_cry_9\
        );

    \I__2388\ : InMux
    port map (
            O => \N__17910\,
            I => \PWMInstance5.un1_periodCounter_2_cry_10\
        );

    \I__2387\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17904\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__17904\,
            I => \N__17901\
        );

    \I__2385\ : Span4Mux_v
    port map (
            O => \N__17901\,
            I => \N__17898\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__17898\,
            I => \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_4\
        );

    \I__2383\ : InMux
    port map (
            O => \N__17895\,
            I => \N__17892\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__17892\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_0\
        );

    \I__2381\ : InMux
    port map (
            O => \N__17889\,
            I => \N__17886\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__17886\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_1\
        );

    \I__2379\ : InMux
    port map (
            O => \N__17883\,
            I => \N__17880\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__17880\,
            I => \N__17877\
        );

    \I__2377\ : Sp12to4
    port map (
            O => \N__17877\,
            I => \N__17874\
        );

    \I__2376\ : Odrv12
    port map (
            O => \N__17874\,
            I => \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_4\
        );

    \I__2375\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17868\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__17868\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_6\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__17865\,
            I => \N__17862\
        );

    \I__2372\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17859\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__17859\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_7\
        );

    \I__2370\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17851\
        );

    \I__2369\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17846\
        );

    \I__2368\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17846\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__17851\,
            I => \PWMInstance5.periodCounterZ0Z_0\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__17846\,
            I => \PWMInstance5.periodCounterZ0Z_0\
        );

    \I__2365\ : InMux
    port map (
            O => \N__17841\,
            I => \PWMInstance5.un1_periodCounter_2_cry_0\
        );

    \I__2364\ : InMux
    port map (
            O => \N__17838\,
            I => \PWMInstance5.un1_periodCounter_2_cry_1\
        );

    \I__2363\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17832\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__17832\,
            I => \N__17829\
        );

    \I__2361\ : Odrv12
    port map (
            O => \N__17829\,
            I => \QuadInstance7.un1_Quad_axb_15\
        );

    \I__2360\ : InMux
    port map (
            O => \N__17826\,
            I => \QuadInstance7.un1_Quad_cry_14\
        );

    \I__2359\ : InMux
    port map (
            O => \N__17823\,
            I => \N__17817\
        );

    \I__2358\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17817\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__17817\,
            I => \pwmWrite_fastZ0Z_1\
        );

    \I__2356\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17808\
        );

    \I__2355\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17808\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__17808\,
            I => \N__17804\
        );

    \I__2353\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17801\
        );

    \I__2352\ : Span4Mux_h
    port map (
            O => \N__17804\,
            I => \N__17798\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__17801\,
            I => \N__17795\
        );

    \I__2350\ : Span4Mux_h
    port map (
            O => \N__17798\,
            I => \N__17792\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__17795\,
            I => \N__17789\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__17792\,
            I => \pwmWriteZ0Z_7\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__17789\,
            I => \pwmWriteZ0Z_7\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__17784\,
            I => \N__17781\
        );

    \I__2345\ : InMux
    port map (
            O => \N__17781\,
            I => \N__17778\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__17778\,
            I => \QuadInstance7.Quad_RNIEBVV2Z0Z_7\
        );

    \I__2343\ : InMux
    port map (
            O => \N__17775\,
            I => \QuadInstance7.un1_Quad_cry_6\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__17772\,
            I => \N__17769\
        );

    \I__2341\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17766\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__17766\,
            I => \QuadInstance7.Quad_RNIFCVV2Z0Z_8\
        );

    \I__2339\ : InMux
    port map (
            O => \N__17763\,
            I => \bfn_9_9_0_\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__17760\,
            I => \N__17757\
        );

    \I__2337\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17754\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__17754\,
            I => \QuadInstance7.Quad_RNIGDVV2Z0Z_9\
        );

    \I__2335\ : InMux
    port map (
            O => \N__17751\,
            I => \QuadInstance7.un1_Quad_cry_8\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__17748\,
            I => \N__17745\
        );

    \I__2333\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17742\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__17742\,
            I => \QuadInstance7.Quad_RNIOIKU2Z0Z_10\
        );

    \I__2331\ : InMux
    port map (
            O => \N__17739\,
            I => \QuadInstance7.un1_Quad_cry_9\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__17736\,
            I => \N__17733\
        );

    \I__2329\ : InMux
    port map (
            O => \N__17733\,
            I => \N__17730\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__17730\,
            I => \QuadInstance7.Quad_RNIPJKU2Z0Z_11\
        );

    \I__2327\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17724\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__17724\,
            I => \N__17721\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__17721\,
            I => \QuadInstance7.Quad_RNO_0_7_11\
        );

    \I__2324\ : InMux
    port map (
            O => \N__17718\,
            I => \QuadInstance7.un1_Quad_cry_10\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__17715\,
            I => \N__17712\
        );

    \I__2322\ : InMux
    port map (
            O => \N__17712\,
            I => \N__17709\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__17709\,
            I => \QuadInstance7.Quad_RNIQKKU2Z0Z_12\
        );

    \I__2320\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17703\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__17703\,
            I => \N__17700\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__17700\,
            I => \QuadInstance7.Quad_RNO_0_7_12\
        );

    \I__2317\ : InMux
    port map (
            O => \N__17697\,
            I => \QuadInstance7.un1_Quad_cry_11\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__17694\,
            I => \N__17691\
        );

    \I__2315\ : InMux
    port map (
            O => \N__17691\,
            I => \N__17688\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__17688\,
            I => \QuadInstance7.Quad_RNIRLKU2Z0Z_13\
        );

    \I__2313\ : InMux
    port map (
            O => \N__17685\,
            I => \QuadInstance7.un1_Quad_cry_12\
        );

    \I__2312\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17679\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__17679\,
            I => \QuadInstance7.Quad_RNISMKU2Z0Z_14\
        );

    \I__2310\ : InMux
    port map (
            O => \N__17676\,
            I => \QuadInstance7.un1_Quad_cry_13\
        );

    \I__2309\ : CascadeMux
    port map (
            O => \N__17673\,
            I => \N__17670\
        );

    \I__2308\ : InMux
    port map (
            O => \N__17670\,
            I => \N__17667\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__17667\,
            I => \QuadInstance7.Quad_RNI85VV2Z0Z_1\
        );

    \I__2306\ : InMux
    port map (
            O => \N__17664\,
            I => \QuadInstance7.un1_Quad_cry_0\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__17661\,
            I => \N__17658\
        );

    \I__2304\ : InMux
    port map (
            O => \N__17658\,
            I => \N__17655\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__17655\,
            I => \QuadInstance7.Quad_RNI96VV2Z0Z_2\
        );

    \I__2302\ : InMux
    port map (
            O => \N__17652\,
            I => \QuadInstance7.un1_Quad_cry_1\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__17649\,
            I => \N__17646\
        );

    \I__2300\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17643\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__17643\,
            I => \QuadInstance7.Quad_RNIA7VV2Z0Z_3\
        );

    \I__2298\ : InMux
    port map (
            O => \N__17640\,
            I => \QuadInstance7.un1_Quad_cry_2\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__17637\,
            I => \N__17634\
        );

    \I__2296\ : InMux
    port map (
            O => \N__17634\,
            I => \N__17631\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__17631\,
            I => \QuadInstance7.Quad_RNIB8VV2Z0Z_4\
        );

    \I__2294\ : InMux
    port map (
            O => \N__17628\,
            I => \QuadInstance7.un1_Quad_cry_3\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__17625\,
            I => \N__17622\
        );

    \I__2292\ : InMux
    port map (
            O => \N__17622\,
            I => \N__17619\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__17619\,
            I => \QuadInstance7.Quad_RNIC9VV2Z0Z_5\
        );

    \I__2290\ : InMux
    port map (
            O => \N__17616\,
            I => \QuadInstance7.un1_Quad_cry_4\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__17613\,
            I => \N__17610\
        );

    \I__2288\ : InMux
    port map (
            O => \N__17610\,
            I => \N__17607\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__17607\,
            I => \QuadInstance7.Quad_RNIDAVV2Z0Z_6\
        );

    \I__2286\ : InMux
    port map (
            O => \N__17604\,
            I => \QuadInstance7.un1_Quad_cry_5\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__17601\,
            I => \N__17598\
        );

    \I__2284\ : InMux
    port map (
            O => \N__17598\,
            I => \N__17595\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__17595\,
            I => \N__17585\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__17594\,
            I => \N__17581\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__17593\,
            I => \N__17578\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__17592\,
            I => \N__17573\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__17591\,
            I => \N__17569\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__17590\,
            I => \N__17565\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__17589\,
            I => \N__17562\
        );

    \I__2276\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17558\
        );

    \I__2275\ : Span4Mux_h
    port map (
            O => \N__17585\,
            I => \N__17555\
        );

    \I__2274\ : InMux
    port map (
            O => \N__17584\,
            I => \N__17546\
        );

    \I__2273\ : InMux
    port map (
            O => \N__17581\,
            I => \N__17546\
        );

    \I__2272\ : InMux
    port map (
            O => \N__17578\,
            I => \N__17546\
        );

    \I__2271\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17546\
        );

    \I__2270\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17529\
        );

    \I__2269\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17529\
        );

    \I__2268\ : InMux
    port map (
            O => \N__17572\,
            I => \N__17529\
        );

    \I__2267\ : InMux
    port map (
            O => \N__17569\,
            I => \N__17529\
        );

    \I__2266\ : InMux
    port map (
            O => \N__17568\,
            I => \N__17529\
        );

    \I__2265\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17529\
        );

    \I__2264\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17529\
        );

    \I__2263\ : InMux
    port map (
            O => \N__17561\,
            I => \N__17529\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__17558\,
            I => \QuadInstance2.un1_count_enable_i_a2_0_1\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__17555\,
            I => \QuadInstance2.un1_count_enable_i_a2_0_1\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__17546\,
            I => \QuadInstance2.un1_count_enable_i_a2_0_1\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__17529\,
            I => \QuadInstance2.un1_count_enable_i_a2_0_1\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__17520\,
            I => \N__17517\
        );

    \I__2257\ : InMux
    port map (
            O => \N__17517\,
            I => \N__17514\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__17514\,
            I => \N__17511\
        );

    \I__2255\ : Span4Mux_h
    port map (
            O => \N__17511\,
            I => \N__17508\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__17508\,
            I => \QuadInstance2.Quad_RNIJ03G2Z0Z_13\
        );

    \I__2253\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17490\
        );

    \I__2252\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17490\
        );

    \I__2251\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17490\
        );

    \I__2250\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17490\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__17501\,
            I => \N__17487\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__17500\,
            I => \N__17483\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__17499\,
            I => \N__17479\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__17490\,
            I => \N__17471\
        );

    \I__2245\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17466\
        );

    \I__2244\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17466\
        );

    \I__2243\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17457\
        );

    \I__2242\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17457\
        );

    \I__2241\ : InMux
    port map (
            O => \N__17479\,
            I => \N__17457\
        );

    \I__2240\ : InMux
    port map (
            O => \N__17478\,
            I => \N__17457\
        );

    \I__2239\ : InMux
    port map (
            O => \N__17477\,
            I => \N__17448\
        );

    \I__2238\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17448\
        );

    \I__2237\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17448\
        );

    \I__2236\ : InMux
    port map (
            O => \N__17474\,
            I => \N__17448\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__17471\,
            I => \QuadInstance5.un1_count_enable_i_a2_0_1\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__17466\,
            I => \QuadInstance5.un1_count_enable_i_a2_0_1\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__17457\,
            I => \QuadInstance5.un1_count_enable_i_a2_0_1\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__17448\,
            I => \QuadInstance5.un1_count_enable_i_a2_0_1\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__17439\,
            I => \QuadInstance5.un1_count_enable_i_a2_0_1_cascade_\
        );

    \I__2230\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17433\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__17433\,
            I => \N__17430\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__17430\,
            I => \N__17427\
        );

    \I__2227\ : Span4Mux_h
    port map (
            O => \N__17427\,
            I => \N__17424\
        );

    \I__2226\ : Span4Mux_h
    port map (
            O => \N__17424\,
            I => \N__17421\
        );

    \I__2225\ : Odrv4
    port map (
            O => \N__17421\,
            I => \ch7_B_c\
        );

    \I__2224\ : InMux
    port map (
            O => \N__17418\,
            I => \N__17415\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__17415\,
            I => \N__17412\
        );

    \I__2222\ : Odrv12
    port map (
            O => \N__17412\,
            I => \QuadInstance7.delayedCh_BZ0Z_0\
        );

    \I__2221\ : IoInMux
    port map (
            O => \N__17409\,
            I => \N__17406\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__17406\,
            I => \PWM0_obufLegalizeSB_DFFNet\
        );

    \I__2219\ : IoInMux
    port map (
            O => \N__17403\,
            I => \N__17400\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__17400\,
            I => \PWM1_obufLegalizeSB_DFFNet\
        );

    \I__2217\ : IoInMux
    port map (
            O => \N__17397\,
            I => \N__17394\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__17394\,
            I => \PWM6_obufLegalizeSB_DFFNet\
        );

    \I__2215\ : IoInMux
    port map (
            O => \N__17391\,
            I => \N__17388\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__17388\,
            I => \PWM7_obufLegalizeSB_DFFNet\
        );

    \I__2213\ : InMux
    port map (
            O => \N__17385\,
            I => \N__17382\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__17382\,
            I => \N__17379\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__17379\,
            I => \ch3_B_c\
        );

    \I__2210\ : InMux
    port map (
            O => \N__17376\,
            I => \N__17373\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__17373\,
            I => \N__17370\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__17370\,
            I => \N__17367\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__17367\,
            I => \QuadInstance2.Quad_RNO_0_2_4\
        );

    \I__2206\ : InMux
    port map (
            O => \N__17364\,
            I => \N__17361\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__17361\,
            I => \N__17358\
        );

    \I__2204\ : Span4Mux_h
    port map (
            O => \N__17358\,
            I => \N__17355\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__17355\,
            I => \ch5_A_c\
        );

    \I__2202\ : InMux
    port map (
            O => \N__17352\,
            I => \N__17349\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__17349\,
            I => \QuadInstance5.delayedCh_AZ0Z_0\
        );

    \I__2200\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17343\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__17343\,
            I => \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNOZ0\
        );

    \I__2198\ : InMux
    port map (
            O => \N__17340\,
            I => \N__17337\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__17337\,
            I => \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNOZ0\
        );

    \I__2196\ : InMux
    port map (
            O => \N__17334\,
            I => \N__17331\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__17331\,
            I => \N__17328\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__17328\,
            I => \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNOZ0\
        );

    \I__2193\ : InMux
    port map (
            O => \N__17325\,
            I => \N__17322\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__17322\,
            I => \N__17319\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__17319\,
            I => \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNOZ0\
        );

    \I__2190\ : InMux
    port map (
            O => \N__17316\,
            I => \N__17313\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__17313\,
            I => \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNOZ0\
        );

    \I__2188\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17307\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__17307\,
            I => \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNOZ0\
        );

    \I__2186\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17301\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__17301\,
            I => \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNOZ0\
        );

    \I__2184\ : InMux
    port map (
            O => \N__17298\,
            I => \N__17295\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__17295\,
            I => \PWMInstance0.un1_periodCounter12_1_0_a2_0\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__17292\,
            I => \N__17285\
        );

    \I__2181\ : InMux
    port map (
            O => \N__17291\,
            I => \N__17281\
        );

    \I__2180\ : InMux
    port map (
            O => \N__17290\,
            I => \N__17278\
        );

    \I__2179\ : InMux
    port map (
            O => \N__17289\,
            I => \N__17273\
        );

    \I__2178\ : InMux
    port map (
            O => \N__17288\,
            I => \N__17273\
        );

    \I__2177\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17270\
        );

    \I__2176\ : InMux
    port map (
            O => \N__17284\,
            I => \N__17267\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__17281\,
            I => \N__17260\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__17278\,
            I => \N__17260\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__17273\,
            I => \N__17260\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__17270\,
            I => \PWMInstance0.out_0_sqmuxa\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__17267\,
            I => \PWMInstance0.out_0_sqmuxa\
        );

    \I__2170\ : Odrv12
    port map (
            O => \N__17260\,
            I => \PWMInstance0.out_0_sqmuxa\
        );

    \I__2169\ : InMux
    port map (
            O => \N__17253\,
            I => \bfn_8_16_0_\
        );

    \I__2168\ : IoInMux
    port map (
            O => \N__17250\,
            I => \N__17247\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__17247\,
            I => \N__17244\
        );

    \I__2166\ : Span4Mux_s2_v
    port map (
            O => \N__17244\,
            I => \N__17240\
        );

    \I__2165\ : InMux
    port map (
            O => \N__17243\,
            I => \N__17237\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__17240\,
            I => \PWM0_c\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__17237\,
            I => \PWM0_c\
        );

    \I__2162\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17229\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__17229\,
            I => \N__17226\
        );

    \I__2160\ : Span4Mux_h
    port map (
            O => \N__17226\,
            I => \N__17223\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__17223\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_12\
        );

    \I__2158\ : InMux
    port map (
            O => \N__17220\,
            I => \N__17217\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__17217\,
            I => \N__17214\
        );

    \I__2156\ : Span12Mux_s4_v
    port map (
            O => \N__17214\,
            I => \N__17211\
        );

    \I__2155\ : Odrv12
    port map (
            O => \N__17211\,
            I => \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_4\
        );

    \I__2154\ : InMux
    port map (
            O => \N__17208\,
            I => \N__17205\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__17205\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_6\
        );

    \I__2152\ : InMux
    port map (
            O => \N__17202\,
            I => \N__17199\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__17199\,
            I => \N__17195\
        );

    \I__2150\ : InMux
    port map (
            O => \N__17198\,
            I => \N__17191\
        );

    \I__2149\ : Span4Mux_h
    port map (
            O => \N__17195\,
            I => \N__17188\
        );

    \I__2148\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17185\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__17191\,
            I => \PWMInstance0.periodCounterZ0Z_7\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__17188\,
            I => \PWMInstance0.periodCounterZ0Z_7\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__17185\,
            I => \PWMInstance0.periodCounterZ0Z_7\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__17178\,
            I => \N__17175\
        );

    \I__2143\ : InMux
    port map (
            O => \N__17175\,
            I => \N__17172\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__17172\,
            I => \N__17167\
        );

    \I__2141\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17164\
        );

    \I__2140\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17161\
        );

    \I__2139\ : Span4Mux_h
    port map (
            O => \N__17167\,
            I => \N__17156\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__17164\,
            I => \N__17156\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__17161\,
            I => \PWMInstance0.periodCounterZ0Z_15\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__17156\,
            I => \PWMInstance0.periodCounterZ0Z_15\
        );

    \I__2135\ : InMux
    port map (
            O => \N__17151\,
            I => \N__17148\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__17148\,
            I => \N__17143\
        );

    \I__2133\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17140\
        );

    \I__2132\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17137\
        );

    \I__2131\ : Span4Mux_h
    port map (
            O => \N__17143\,
            I => \N__17134\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__17140\,
            I => \N__17131\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__17137\,
            I => \PWMInstance0.periodCounterZ0Z_14\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__17134\,
            I => \PWMInstance0.periodCounterZ0Z_14\
        );

    \I__2127\ : Odrv12
    port map (
            O => \N__17131\,
            I => \PWMInstance0.periodCounterZ0Z_14\
        );

    \I__2126\ : InMux
    port map (
            O => \N__17124\,
            I => \N__17121\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__17121\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_14\
        );

    \I__2124\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17115\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__17115\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_15\
        );

    \I__2122\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17107\
        );

    \I__2121\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17104\
        );

    \I__2120\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17101\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__17107\,
            I => \N__17098\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__17104\,
            I => \N__17095\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__17101\,
            I => \PWMInstance0.periodCounterZ0Z_10\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__17098\,
            I => \PWMInstance0.periodCounterZ0Z_10\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__17095\,
            I => \PWMInstance0.periodCounterZ0Z_10\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__17088\,
            I => \N__17084\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__17087\,
            I => \N__17081\
        );

    \I__2112\ : InMux
    port map (
            O => \N__17084\,
            I => \N__17077\
        );

    \I__2111\ : InMux
    port map (
            O => \N__17081\,
            I => \N__17074\
        );

    \I__2110\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17071\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__17077\,
            I => \N__17068\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__17074\,
            I => \N__17065\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__17071\,
            I => \PWMInstance0.periodCounterZ0Z_11\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__17068\,
            I => \PWMInstance0.periodCounterZ0Z_11\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__17065\,
            I => \PWMInstance0.periodCounterZ0Z_11\
        );

    \I__2104\ : InMux
    port map (
            O => \N__17058\,
            I => \N__17055\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__17055\,
            I => \N__17052\
        );

    \I__2102\ : Span4Mux_h
    port map (
            O => \N__17052\,
            I => \N__17049\
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__17049\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_10\
        );

    \I__2100\ : InMux
    port map (
            O => \N__17046\,
            I => \N__17043\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__17043\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_11\
        );

    \I__2098\ : InMux
    port map (
            O => \N__17040\,
            I => \N__17037\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__17037\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_13\
        );

    \I__2096\ : InMux
    port map (
            O => \N__17034\,
            I => \N__17031\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__17031\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_12\
        );

    \I__2094\ : InMux
    port map (
            O => \N__17028\,
            I => \N__17023\
        );

    \I__2093\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17020\
        );

    \I__2092\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17017\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__17023\,
            I => \N__17014\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__17020\,
            I => \N__17011\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__17017\,
            I => \PWMInstance0.periodCounterZ0Z_12\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__17014\,
            I => \PWMInstance0.periodCounterZ0Z_12\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__17011\,
            I => \PWMInstance0.periodCounterZ0Z_12\
        );

    \I__2086\ : InMux
    port map (
            O => \N__17004\,
            I => \N__16996\
        );

    \I__2085\ : InMux
    port map (
            O => \N__17003\,
            I => \N__16991\
        );

    \I__2084\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16991\
        );

    \I__2083\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16988\
        );

    \I__2082\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16985\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__16999\,
            I => \N__16982\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__16996\,
            I => \N__16973\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__16991\,
            I => \N__16973\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__16988\,
            I => \N__16973\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__16985\,
            I => \N__16973\
        );

    \I__2076\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16970\
        );

    \I__2075\ : Span12Mux_s5_v
    port map (
            O => \N__16973\,
            I => \N__16967\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__16970\,
            I => \PWMInstance1.out_0_sqmuxa\
        );

    \I__2073\ : Odrv12
    port map (
            O => \N__16967\,
            I => \PWMInstance1.out_0_sqmuxa\
        );

    \I__2072\ : InMux
    port map (
            O => \N__16962\,
            I => \N__16959\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__16959\,
            I => \N__16956\
        );

    \I__2070\ : Odrv12
    port map (
            O => \N__16956\,
            I => \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_4\
        );

    \I__2069\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16950\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__16950\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_2\
        );

    \I__2067\ : InMux
    port map (
            O => \N__16947\,
            I => \N__16944\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__16944\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_3\
        );

    \I__2065\ : InMux
    port map (
            O => \N__16941\,
            I => \N__16938\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__16938\,
            I => \N__16935\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__16935\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_14\
        );

    \I__2062\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16929\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__16929\,
            I => \N__16926\
        );

    \I__2060\ : Span12Mux_s3_v
    port map (
            O => \N__16926\,
            I => \N__16923\
        );

    \I__2059\ : Odrv12
    port map (
            O => \N__16923\,
            I => \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_4\
        );

    \I__2058\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16917\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__16917\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_15\
        );

    \I__2056\ : InMux
    port map (
            O => \N__16914\,
            I => \N__16911\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__16911\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_9\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__16908\,
            I => \N__16905\
        );

    \I__2053\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16901\
        );

    \I__2052\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16897\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__16901\,
            I => \N__16894\
        );

    \I__2050\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16891\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__16897\,
            I => \N__16886\
        );

    \I__2048\ : Span4Mux_h
    port map (
            O => \N__16894\,
            I => \N__16886\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__16891\,
            I => \PWMInstance0.periodCounterZ0Z_9\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__16886\,
            I => \PWMInstance0.periodCounterZ0Z_9\
        );

    \I__2045\ : InMux
    port map (
            O => \N__16881\,
            I => \N__16878\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__16878\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_8\
        );

    \I__2043\ : InMux
    port map (
            O => \N__16875\,
            I => \N__16869\
        );

    \I__2042\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16869\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__16869\,
            I => \N__16866\
        );

    \I__2040\ : Span4Mux_h
    port map (
            O => \N__16866\,
            I => \N__16862\
        );

    \I__2039\ : InMux
    port map (
            O => \N__16865\,
            I => \N__16859\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__16862\,
            I => \pwmWriteZ0Z_0\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__16859\,
            I => \pwmWriteZ0Z_0\
        );

    \I__2036\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16850\
        );

    \I__2035\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16847\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__16850\,
            I => \QuadInstance7.delayedCh_BZ0Z_1\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__16847\,
            I => \QuadInstance7.delayedCh_BZ0Z_1\
        );

    \I__2032\ : InMux
    port map (
            O => \N__16842\,
            I => \N__16836\
        );

    \I__2031\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16836\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__16836\,
            I => \QuadInstance7.delayedCh_BZ0Z_2\
        );

    \I__2029\ : InMux
    port map (
            O => \N__16833\,
            I => \N__16830\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__16830\,
            I => \PWMInstance1.un1_periodCounter12_1_0_a2_0\
        );

    \I__2027\ : CEMux
    port map (
            O => \N__16827\,
            I => \N__16819\
        );

    \I__2026\ : CEMux
    port map (
            O => \N__16826\,
            I => \N__16816\
        );

    \I__2025\ : CEMux
    port map (
            O => \N__16825\,
            I => \N__16813\
        );

    \I__2024\ : CEMux
    port map (
            O => \N__16824\,
            I => \N__16810\
        );

    \I__2023\ : CEMux
    port map (
            O => \N__16823\,
            I => \N__16807\
        );

    \I__2022\ : CEMux
    port map (
            O => \N__16822\,
            I => \N__16804\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__16819\,
            I => \N__16800\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__16816\,
            I => \N__16795\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__16813\,
            I => \N__16795\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__16810\,
            I => \N__16792\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__16807\,
            I => \N__16789\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__16804\,
            I => \N__16786\
        );

    \I__2015\ : CEMux
    port map (
            O => \N__16803\,
            I => \N__16783\
        );

    \I__2014\ : Span4Mux_s3_v
    port map (
            O => \N__16800\,
            I => \N__16778\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__16795\,
            I => \N__16778\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__16792\,
            I => \N__16775\
        );

    \I__2011\ : Span4Mux_s2_v
    port map (
            O => \N__16789\,
            I => \N__16768\
        );

    \I__2010\ : Span4Mux_h
    port map (
            O => \N__16786\,
            I => \N__16768\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__16783\,
            I => \N__16768\
        );

    \I__2008\ : Span4Mux_v
    port map (
            O => \N__16778\,
            I => \N__16765\
        );

    \I__2007\ : Span4Mux_h
    port map (
            O => \N__16775\,
            I => \N__16760\
        );

    \I__2006\ : Span4Mux_v
    port map (
            O => \N__16768\,
            I => \N__16760\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__16765\,
            I => \PWMInstance1.pwmWrite_0_1\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__16760\,
            I => \PWMInstance1.pwmWrite_0_1\
        );

    \I__2003\ : InMux
    port map (
            O => \N__16755\,
            I => \N__16746\
        );

    \I__2002\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16746\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16746\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__16746\,
            I => \pwmWriteZ0Z_1\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__16743\,
            I => \N__16739\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__16742\,
            I => \N__16736\
        );

    \I__1997\ : InMux
    port map (
            O => \N__16739\,
            I => \N__16725\
        );

    \I__1996\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16725\
        );

    \I__1995\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16725\
        );

    \I__1994\ : InMux
    port map (
            O => \N__16734\,
            I => \N__16725\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__16725\,
            I => \PWMInstance1.clkCountZ0Z_1\
        );

    \I__1992\ : InMux
    port map (
            O => \N__16722\,
            I => \N__16710\
        );

    \I__1991\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16710\
        );

    \I__1990\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16710\
        );

    \I__1989\ : InMux
    port map (
            O => \N__16719\,
            I => \N__16710\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__16710\,
            I => \PWMInstance1.clkCountZ0Z_0\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__16707\,
            I => \N__16704\
        );

    \I__1986\ : InMux
    port map (
            O => \N__16704\,
            I => \N__16697\
        );

    \I__1985\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16697\
        );

    \I__1984\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16694\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__16697\,
            I => \N__16691\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__16694\,
            I => \PWMInstance1.periodCounterZ0Z_16\
        );

    \I__1981\ : Odrv12
    port map (
            O => \N__16691\,
            I => \PWMInstance1.periodCounterZ0Z_16\
        );

    \I__1980\ : InMux
    port map (
            O => \N__16686\,
            I => \N__16683\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__16683\,
            I => \N__16679\
        );

    \I__1978\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16675\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__16679\,
            I => \N__16672\
        );

    \I__1976\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16669\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__16675\,
            I => \N__16664\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__16672\,
            I => \N__16664\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__16669\,
            I => \PWMInstance1.periodCounterZ0Z_7\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__16664\,
            I => \PWMInstance1.periodCounterZ0Z_7\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__16659\,
            I => \N__16656\
        );

    \I__1970\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16652\
        );

    \I__1969\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16649\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__16652\,
            I => \N__16645\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__16649\,
            I => \N__16642\
        );

    \I__1966\ : InMux
    port map (
            O => \N__16648\,
            I => \N__16639\
        );

    \I__1965\ : Span4Mux_h
    port map (
            O => \N__16645\,
            I => \N__16636\
        );

    \I__1964\ : Span12Mux_s11_v
    port map (
            O => \N__16642\,
            I => \N__16633\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__16639\,
            I => \PWMInstance1.periodCounterZ0Z_15\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__16636\,
            I => \PWMInstance1.periodCounterZ0Z_15\
        );

    \I__1961\ : Odrv12
    port map (
            O => \N__16633\,
            I => \PWMInstance1.periodCounterZ0Z_15\
        );

    \I__1960\ : InMux
    port map (
            O => \N__16626\,
            I => \N__16623\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__16623\,
            I => \N__16620\
        );

    \I__1958\ : Span4Mux_v
    port map (
            O => \N__16620\,
            I => \N__16615\
        );

    \I__1957\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16612\
        );

    \I__1956\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16609\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__16615\,
            I => \N__16604\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__16612\,
            I => \N__16604\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__16609\,
            I => \PWMInstance1.periodCounterZ0Z_1\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__16604\,
            I => \PWMInstance1.periodCounterZ0Z_1\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__16599\,
            I => \PWMInstance1.un1_periodCounter12_1_0_a2_0_6_cascade_\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__16596\,
            I => \N__16592\
        );

    \I__1949\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16589\
        );

    \I__1948\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16586\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__16589\,
            I => \N__16581\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__16586\,
            I => \N__16581\
        );

    \I__1945\ : Span12Mux_s2_v
    port map (
            O => \N__16581\,
            I => \N__16577\
        );

    \I__1944\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16574\
        );

    \I__1943\ : Odrv12
    port map (
            O => \N__16577\,
            I => \PWMInstance1.periodCounter12\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__16574\,
            I => \PWMInstance1.periodCounter12\
        );

    \I__1941\ : InMux
    port map (
            O => \N__16569\,
            I => \N__16566\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__16566\,
            I => \N__16563\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__16563\,
            I => \N__16560\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__16560\,
            I => \N__16557\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__16557\,
            I => \PWMInstance1.un1_periodCounter12_1_0_a2_0_10\
        );

    \I__1936\ : InMux
    port map (
            O => \N__16554\,
            I => \N__16551\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__16551\,
            I => \N__16548\
        );

    \I__1934\ : Span12Mux_h
    port map (
            O => \N__16548\,
            I => \N__16545\
        );

    \I__1933\ : Odrv12
    port map (
            O => \N__16545\,
            I => \PWMInstance1.un1_periodCounter12_1_0_a2_0_9\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__16542\,
            I => \PWMInstance1.un1_periodCounter12_1_0_a2_0_14_cascade_\
        );

    \I__1931\ : InMux
    port map (
            O => \N__16539\,
            I => \N__16536\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__16536\,
            I => \N__16533\
        );

    \I__1929\ : Span4Mux_v
    port map (
            O => \N__16533\,
            I => \N__16530\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__16530\,
            I => \N__16527\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__16527\,
            I => \PWMInstance1.un1_periodCounter12_1_0_a2_0_12\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__16524\,
            I => \N__16518\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__16523\,
            I => \N__16515\
        );

    \I__1924\ : InMux
    port map (
            O => \N__16522\,
            I => \N__16502\
        );

    \I__1923\ : InMux
    port map (
            O => \N__16521\,
            I => \N__16495\
        );

    \I__1922\ : InMux
    port map (
            O => \N__16518\,
            I => \N__16495\
        );

    \I__1921\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16495\
        );

    \I__1920\ : InMux
    port map (
            O => \N__16514\,
            I => \N__16484\
        );

    \I__1919\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16484\
        );

    \I__1918\ : InMux
    port map (
            O => \N__16512\,
            I => \N__16484\
        );

    \I__1917\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16484\
        );

    \I__1916\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16484\
        );

    \I__1915\ : InMux
    port map (
            O => \N__16509\,
            I => \N__16473\
        );

    \I__1914\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16473\
        );

    \I__1913\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16473\
        );

    \I__1912\ : InMux
    port map (
            O => \N__16506\,
            I => \N__16473\
        );

    \I__1911\ : InMux
    port map (
            O => \N__16505\,
            I => \N__16473\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__16502\,
            I => \QuadInstance7.un1_count_enable_i_a2_0_1\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__16495\,
            I => \QuadInstance7.un1_count_enable_i_a2_0_1\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__16484\,
            I => \QuadInstance7.un1_count_enable_i_a2_0_1\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__16473\,
            I => \QuadInstance7.un1_count_enable_i_a2_0_1\
        );

    \I__1906\ : InMux
    port map (
            O => \N__16464\,
            I => \N__16459\
        );

    \I__1905\ : InMux
    port map (
            O => \N__16463\,
            I => \N__16454\
        );

    \I__1904\ : InMux
    port map (
            O => \N__16462\,
            I => \N__16454\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__16459\,
            I => \QuadInstance7.delayedCh_AZ0Z_1\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__16454\,
            I => \QuadInstance7.delayedCh_AZ0Z_1\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__16449\,
            I => \N__16446\
        );

    \I__1900\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16443\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__16443\,
            I => \QuadInstance7.delayedCh_AZ0Z_2\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__16440\,
            I => \QuadInstance7.un1_count_enable_i_a2_0_1_cascade_\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__16437\,
            I => \QuadInstance7.count_enable_cascade_\
        );

    \I__1896\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16431\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__16431\,
            I => \QuadInstance2.Quad_RNO_0_2_10\
        );

    \I__1894\ : InMux
    port map (
            O => \N__16428\,
            I => \N__16425\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__16425\,
            I => \QuadInstance2.Quad_RNO_0_2_14\
        );

    \I__1892\ : InMux
    port map (
            O => \N__16422\,
            I => \N__16419\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__16419\,
            I => \QuadInstance2.Quad_RNO_0_2_12\
        );

    \I__1890\ : InMux
    port map (
            O => \N__16416\,
            I => \N__16413\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__16413\,
            I => \N__16410\
        );

    \I__1888\ : Span12Mux_h
    port map (
            O => \N__16410\,
            I => \N__16407\
        );

    \I__1887\ : Odrv12
    port map (
            O => \N__16407\,
            I => \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_4\
        );

    \I__1886\ : InMux
    port map (
            O => \N__16404\,
            I => \bfn_8_5_0_\
        );

    \I__1885\ : IoInMux
    port map (
            O => \N__16401\,
            I => \N__16398\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__16398\,
            I => \N__16395\
        );

    \I__1883\ : Span4Mux_s3_v
    port map (
            O => \N__16395\,
            I => \N__16392\
        );

    \I__1882\ : Sp12to4
    port map (
            O => \N__16392\,
            I => \N__16389\
        );

    \I__1881\ : Span12Mux_h
    port map (
            O => \N__16389\,
            I => \N__16386\
        );

    \I__1880\ : Span12Mux_v
    port map (
            O => \N__16386\,
            I => \N__16382\
        );

    \I__1879\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16379\
        );

    \I__1878\ : Odrv12
    port map (
            O => \N__16382\,
            I => \PWM5_c\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__16379\,
            I => \PWM5_c\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__16374\,
            I => \N__16371\
        );

    \I__1875\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16368\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__16368\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_12\
        );

    \I__1873\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16362\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__16362\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_10\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__16359\,
            I => \N__16356\
        );

    \I__1870\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16353\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__16353\,
            I => \QuadInstance2.Quad_RNO_0_2_9\
        );

    \I__1868\ : InMux
    port map (
            O => \N__16350\,
            I => \N__16345\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__16349\,
            I => \N__16342\
        );

    \I__1866\ : InMux
    port map (
            O => \N__16348\,
            I => \N__16339\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__16345\,
            I => \N__16336\
        );

    \I__1864\ : InMux
    port map (
            O => \N__16342\,
            I => \N__16333\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__16339\,
            I => \PWMInstance1.periodCounterZ0Z_11\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__16336\,
            I => \PWMInstance1.periodCounterZ0Z_11\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__16333\,
            I => \PWMInstance1.periodCounterZ0Z_11\
        );

    \I__1860\ : InMux
    port map (
            O => \N__16326\,
            I => \PWMInstance1.un1_periodCounter_2_cry_10\
        );

    \I__1859\ : InMux
    port map (
            O => \N__16323\,
            I => \N__16319\
        );

    \I__1858\ : InMux
    port map (
            O => \N__16322\,
            I => \N__16315\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__16319\,
            I => \N__16312\
        );

    \I__1856\ : InMux
    port map (
            O => \N__16318\,
            I => \N__16309\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__16315\,
            I => \PWMInstance1.periodCounterZ0Z_12\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__16312\,
            I => \PWMInstance1.periodCounterZ0Z_12\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__16309\,
            I => \PWMInstance1.periodCounterZ0Z_12\
        );

    \I__1852\ : InMux
    port map (
            O => \N__16302\,
            I => \PWMInstance1.un1_periodCounter_2_cry_11\
        );

    \I__1851\ : InMux
    port map (
            O => \N__16299\,
            I => \N__16296\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__16296\,
            I => \N__16291\
        );

    \I__1849\ : InMux
    port map (
            O => \N__16295\,
            I => \N__16288\
        );

    \I__1848\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16285\
        );

    \I__1847\ : Span4Mux_h
    port map (
            O => \N__16291\,
            I => \N__16280\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__16288\,
            I => \N__16280\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__16285\,
            I => \PWMInstance1.periodCounterZ0Z_13\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__16280\,
            I => \PWMInstance1.periodCounterZ0Z_13\
        );

    \I__1843\ : InMux
    port map (
            O => \N__16275\,
            I => \PWMInstance1.un1_periodCounter_2_cry_12\
        );

    \I__1842\ : InMux
    port map (
            O => \N__16272\,
            I => \N__16268\
        );

    \I__1841\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16264\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__16268\,
            I => \N__16261\
        );

    \I__1839\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16258\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__16264\,
            I => \PWMInstance1.periodCounterZ0Z_14\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__16261\,
            I => \PWMInstance1.periodCounterZ0Z_14\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__16258\,
            I => \PWMInstance1.periodCounterZ0Z_14\
        );

    \I__1835\ : InMux
    port map (
            O => \N__16251\,
            I => \PWMInstance1.un1_periodCounter_2_cry_13\
        );

    \I__1834\ : InMux
    port map (
            O => \N__16248\,
            I => \PWMInstance1.un1_periodCounter_2_cry_14\
        );

    \I__1833\ : InMux
    port map (
            O => \N__16245\,
            I => \bfn_8_3_0_\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__16242\,
            I => \N__16237\
        );

    \I__1831\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16234\
        );

    \I__1830\ : InMux
    port map (
            O => \N__16240\,
            I => \N__16229\
        );

    \I__1829\ : InMux
    port map (
            O => \N__16237\,
            I => \N__16229\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__16234\,
            I => \PWMInstance1.periodCounterZ0Z_3\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__16229\,
            I => \PWMInstance1.periodCounterZ0Z_3\
        );

    \I__1826\ : InMux
    port map (
            O => \N__16224\,
            I => \PWMInstance1.un1_periodCounter_2_cry_2\
        );

    \I__1825\ : InMux
    port map (
            O => \N__16221\,
            I => \N__16216\
        );

    \I__1824\ : InMux
    port map (
            O => \N__16220\,
            I => \N__16211\
        );

    \I__1823\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16211\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__16216\,
            I => \PWMInstance1.periodCounterZ0Z_4\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__16211\,
            I => \PWMInstance1.periodCounterZ0Z_4\
        );

    \I__1820\ : InMux
    port map (
            O => \N__16206\,
            I => \PWMInstance1.un1_periodCounter_2_cry_3\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__16203\,
            I => \N__16198\
        );

    \I__1818\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16195\
        );

    \I__1817\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16190\
        );

    \I__1816\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16190\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__16195\,
            I => \PWMInstance1.periodCounterZ0Z_5\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__16190\,
            I => \PWMInstance1.periodCounterZ0Z_5\
        );

    \I__1813\ : InMux
    port map (
            O => \N__16185\,
            I => \PWMInstance1.un1_periodCounter_2_cry_4\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__16182\,
            I => \N__16179\
        );

    \I__1811\ : InMux
    port map (
            O => \N__16179\,
            I => \N__16173\
        );

    \I__1810\ : InMux
    port map (
            O => \N__16178\,
            I => \N__16173\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__16173\,
            I => \N__16169\
        );

    \I__1808\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16166\
        );

    \I__1807\ : Span4Mux_h
    port map (
            O => \N__16169\,
            I => \N__16163\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__16166\,
            I => \PWMInstance1.periodCounterZ0Z_6\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__16163\,
            I => \PWMInstance1.periodCounterZ0Z_6\
        );

    \I__1804\ : InMux
    port map (
            O => \N__16158\,
            I => \PWMInstance1.un1_periodCounter_2_cry_5\
        );

    \I__1803\ : InMux
    port map (
            O => \N__16155\,
            I => \PWMInstance1.un1_periodCounter_2_cry_6\
        );

    \I__1802\ : InMux
    port map (
            O => \N__16152\,
            I => \N__16147\
        );

    \I__1801\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16144\
        );

    \I__1800\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16141\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__16147\,
            I => \PWMInstance1.periodCounterZ0Z_8\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__16144\,
            I => \PWMInstance1.periodCounterZ0Z_8\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__16141\,
            I => \PWMInstance1.periodCounterZ0Z_8\
        );

    \I__1796\ : InMux
    port map (
            O => \N__16134\,
            I => \bfn_8_2_0_\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__16131\,
            I => \N__16126\
        );

    \I__1794\ : InMux
    port map (
            O => \N__16130\,
            I => \N__16123\
        );

    \I__1793\ : InMux
    port map (
            O => \N__16129\,
            I => \N__16120\
        );

    \I__1792\ : InMux
    port map (
            O => \N__16126\,
            I => \N__16117\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__16123\,
            I => \PWMInstance1.periodCounterZ0Z_9\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__16120\,
            I => \PWMInstance1.periodCounterZ0Z_9\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__16117\,
            I => \PWMInstance1.periodCounterZ0Z_9\
        );

    \I__1788\ : InMux
    port map (
            O => \N__16110\,
            I => \PWMInstance1.un1_periodCounter_2_cry_8\
        );

    \I__1787\ : InMux
    port map (
            O => \N__16107\,
            I => \N__16104\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__16104\,
            I => \N__16099\
        );

    \I__1785\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16096\
        );

    \I__1784\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16093\
        );

    \I__1783\ : Span4Mux_h
    port map (
            O => \N__16099\,
            I => \N__16090\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__16096\,
            I => \PWMInstance1.periodCounterZ0Z_10\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__16093\,
            I => \PWMInstance1.periodCounterZ0Z_10\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__16090\,
            I => \PWMInstance1.periodCounterZ0Z_10\
        );

    \I__1779\ : InMux
    port map (
            O => \N__16083\,
            I => \PWMInstance1.un1_periodCounter_2_cry_9\
        );

    \I__1778\ : InMux
    port map (
            O => \N__16080\,
            I => \PWMInstance0.un1_periodCounter_2_cry_10\
        );

    \I__1777\ : InMux
    port map (
            O => \N__16077\,
            I => \PWMInstance0.un1_periodCounter_2_cry_11\
        );

    \I__1776\ : InMux
    port map (
            O => \N__16074\,
            I => \PWMInstance0.un1_periodCounter_2_cry_12\
        );

    \I__1775\ : InMux
    port map (
            O => \N__16071\,
            I => \PWMInstance0.un1_periodCounter_2_cry_13\
        );

    \I__1774\ : InMux
    port map (
            O => \N__16068\,
            I => \PWMInstance0.un1_periodCounter_2_cry_14\
        );

    \I__1773\ : InMux
    port map (
            O => \N__16065\,
            I => \bfn_7_18_0_\
        );

    \I__1772\ : InMux
    port map (
            O => \N__16062\,
            I => \N__16055\
        );

    \I__1771\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16055\
        );

    \I__1770\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16052\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__16055\,
            I => \N__16049\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__16052\,
            I => \PWMInstance0.periodCounterZ0Z_16\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__16049\,
            I => \PWMInstance0.periodCounterZ0Z_16\
        );

    \I__1766\ : InMux
    port map (
            O => \N__16044\,
            I => \N__16037\
        );

    \I__1765\ : InMux
    port map (
            O => \N__16043\,
            I => \N__16037\
        );

    \I__1764\ : InMux
    port map (
            O => \N__16042\,
            I => \N__16034\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__16037\,
            I => \N__16031\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__16034\,
            I => \PWMInstance1.periodCounterZ0Z_0\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__16031\,
            I => \PWMInstance1.periodCounterZ0Z_0\
        );

    \I__1760\ : InMux
    port map (
            O => \N__16026\,
            I => \PWMInstance1.un1_periodCounter_2_cry_0\
        );

    \I__1759\ : InMux
    port map (
            O => \N__16023\,
            I => \N__16018\
        );

    \I__1758\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16013\
        );

    \I__1757\ : InMux
    port map (
            O => \N__16021\,
            I => \N__16013\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__16018\,
            I => \PWMInstance1.periodCounterZ0Z_2\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__16013\,
            I => \PWMInstance1.periodCounterZ0Z_2\
        );

    \I__1754\ : InMux
    port map (
            O => \N__16008\,
            I => \PWMInstance1.un1_periodCounter_2_cry_1\
        );

    \I__1753\ : InMux
    port map (
            O => \N__16005\,
            I => \N__15998\
        );

    \I__1752\ : InMux
    port map (
            O => \N__16004\,
            I => \N__15998\
        );

    \I__1751\ : InMux
    port map (
            O => \N__16003\,
            I => \N__15995\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__15998\,
            I => \N__15992\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__15995\,
            I => \PWMInstance0.periodCounterZ0Z_2\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__15992\,
            I => \PWMInstance0.periodCounterZ0Z_2\
        );

    \I__1747\ : InMux
    port map (
            O => \N__15987\,
            I => \PWMInstance0.un1_periodCounter_2_cry_1\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__15984\,
            I => \N__15980\
        );

    \I__1745\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15974\
        );

    \I__1744\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15974\
        );

    \I__1743\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15971\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__15974\,
            I => \N__15968\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__15971\,
            I => \PWMInstance0.periodCounterZ0Z_3\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__15968\,
            I => \PWMInstance0.periodCounterZ0Z_3\
        );

    \I__1739\ : InMux
    port map (
            O => \N__15963\,
            I => \PWMInstance0.un1_periodCounter_2_cry_2\
        );

    \I__1738\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15953\
        );

    \I__1737\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15953\
        );

    \I__1736\ : InMux
    port map (
            O => \N__15958\,
            I => \N__15950\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__15953\,
            I => \N__15947\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__15950\,
            I => \PWMInstance0.periodCounterZ0Z_4\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__15947\,
            I => \PWMInstance0.periodCounterZ0Z_4\
        );

    \I__1732\ : InMux
    port map (
            O => \N__15942\,
            I => \PWMInstance0.un1_periodCounter_2_cry_3\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__15939\,
            I => \N__15935\
        );

    \I__1730\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15929\
        );

    \I__1729\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15929\
        );

    \I__1728\ : InMux
    port map (
            O => \N__15934\,
            I => \N__15926\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__15929\,
            I => \N__15923\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__15926\,
            I => \PWMInstance0.periodCounterZ0Z_5\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__15923\,
            I => \PWMInstance0.periodCounterZ0Z_5\
        );

    \I__1724\ : InMux
    port map (
            O => \N__15918\,
            I => \PWMInstance0.un1_periodCounter_2_cry_4\
        );

    \I__1723\ : InMux
    port map (
            O => \N__15915\,
            I => \PWMInstance0.un1_periodCounter_2_cry_5\
        );

    \I__1722\ : InMux
    port map (
            O => \N__15912\,
            I => \PWMInstance0.un1_periodCounter_2_cry_6\
        );

    \I__1721\ : InMux
    port map (
            O => \N__15909\,
            I => \bfn_7_17_0_\
        );

    \I__1720\ : InMux
    port map (
            O => \N__15906\,
            I => \PWMInstance0.un1_periodCounter_2_cry_8\
        );

    \I__1719\ : InMux
    port map (
            O => \N__15903\,
            I => \PWMInstance0.un1_periodCounter_2_cry_9\
        );

    \I__1718\ : InMux
    port map (
            O => \N__15900\,
            I => \N__15894\
        );

    \I__1717\ : InMux
    port map (
            O => \N__15899\,
            I => \N__15894\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__15894\,
            I => \N__15891\
        );

    \I__1715\ : Odrv12
    port map (
            O => \N__15891\,
            I => \pwmWrite_fastZ0Z_0\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__15888\,
            I => \N__15883\
        );

    \I__1713\ : InMux
    port map (
            O => \N__15887\,
            I => \N__15873\
        );

    \I__1712\ : InMux
    port map (
            O => \N__15886\,
            I => \N__15873\
        );

    \I__1711\ : InMux
    port map (
            O => \N__15883\,
            I => \N__15873\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15873\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__15873\,
            I => \PWMInstance0.clkCountZ0Z_1\
        );

    \I__1708\ : InMux
    port map (
            O => \N__15870\,
            I => \N__15858\
        );

    \I__1707\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15858\
        );

    \I__1706\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15858\
        );

    \I__1705\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15858\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__15858\,
            I => \PWMInstance0.clkCountZ0Z_0\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__15855\,
            I => \PWMInstance0.periodCounter12_cascade_\
        );

    \I__1702\ : InMux
    port map (
            O => \N__15852\,
            I => \N__15849\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__15849\,
            I => \PWMInstance0.un1_periodCounter12_1_0_a2_0_6\
        );

    \I__1700\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15843\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__15843\,
            I => \PWMInstance0.un1_periodCounter12_1_0_a2_0_10\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__15840\,
            I => \PWMInstance0.un1_periodCounter12_1_0_a2_0_14_cascade_\
        );

    \I__1697\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15834\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__15834\,
            I => \PWMInstance0.un1_periodCounter12_1_0_a2_0_12\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__15831\,
            I => \N__15827\
        );

    \I__1694\ : InMux
    port map (
            O => \N__15830\,
            I => \N__15824\
        );

    \I__1693\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15821\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__15824\,
            I => \PWMInstance0.periodCounter12\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__15821\,
            I => \PWMInstance0.periodCounter12\
        );

    \I__1690\ : InMux
    port map (
            O => \N__15816\,
            I => \PWMInstance0.un1_periodCounter_2_cry_0\
        );

    \I__1689\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15810\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__15810\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_2\
        );

    \I__1687\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15804\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__15804\,
            I => \N__15801\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__15801\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_3\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__15798\,
            I => \PWMInstance0.un1_periodCounter12_1_0_a2_0_0_cascade_\
        );

    \I__1683\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15792\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__15792\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_5\
        );

    \I__1681\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15786\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__15786\,
            I => \PWMInstance0.PWMPulseWidthCountZ0Z_4\
        );

    \I__1679\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15780\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__15780\,
            I => \N__15777\
        );

    \I__1677\ : Sp12to4
    port map (
            O => \N__15777\,
            I => \N__15774\
        );

    \I__1676\ : Odrv12
    port map (
            O => \N__15774\,
            I => \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_0\
        );

    \I__1675\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15768\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__15768\,
            I => \N__15765\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__15765\,
            I => \N__15762\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__15762\,
            I => \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_0\
        );

    \I__1671\ : InMux
    port map (
            O => \N__15759\,
            I => \N__15756\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__15756\,
            I => \N__15753\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__15753\,
            I => \N__15750\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__15750\,
            I => \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_0\
        );

    \I__1667\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15744\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__15744\,
            I => \N__15741\
        );

    \I__1665\ : Odrv12
    port map (
            O => \N__15741\,
            I => \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_0\
        );

    \I__1664\ : InMux
    port map (
            O => \N__15738\,
            I => \bfn_7_12_0_\
        );

    \I__1663\ : IoInMux
    port map (
            O => \N__15735\,
            I => \N__15732\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__15732\,
            I => \N__15729\
        );

    \I__1661\ : Span4Mux_s2_v
    port map (
            O => \N__15729\,
            I => \N__15726\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__15726\,
            I => \N__15722\
        );

    \I__1659\ : InMux
    port map (
            O => \N__15725\,
            I => \N__15719\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__15722\,
            I => \PWM1_c\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__15719\,
            I => \PWM1_c\
        );

    \I__1656\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15711\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__15711\,
            I => \N__15708\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__15708\,
            I => \QuadInstance2.Quad_RNIK13G2Z0Z_14\
        );

    \I__1653\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15701\
        );

    \I__1652\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15698\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__15701\,
            I => \QuadInstance2.delayedCh_BZ0Z_1\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__15698\,
            I => \QuadInstance2.delayedCh_BZ0Z_1\
        );

    \I__1649\ : InMux
    port map (
            O => \N__15693\,
            I => \N__15687\
        );

    \I__1648\ : InMux
    port map (
            O => \N__15692\,
            I => \N__15687\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__15687\,
            I => \QuadInstance2.delayedCh_BZ0Z_2\
        );

    \I__1646\ : InMux
    port map (
            O => \N__15684\,
            I => \N__15681\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__15681\,
            I => \N__15678\
        );

    \I__1644\ : Odrv12
    port map (
            O => \N__15678\,
            I => \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_0\
        );

    \I__1643\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15672\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__15672\,
            I => \N__15669\
        );

    \I__1641\ : Odrv12
    port map (
            O => \N__15669\,
            I => \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_0\
        );

    \I__1640\ : InMux
    port map (
            O => \N__15666\,
            I => \N__15663\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__15663\,
            I => \N__15660\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__15660\,
            I => \N__15657\
        );

    \I__1637\ : Span4Mux_v
    port map (
            O => \N__15657\,
            I => \N__15654\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__15654\,
            I => \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_0\
        );

    \I__1635\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15648\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__15648\,
            I => \N__15645\
        );

    \I__1633\ : Span12Mux_v
    port map (
            O => \N__15645\,
            I => \N__15642\
        );

    \I__1632\ : Odrv12
    port map (
            O => \N__15642\,
            I => \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_0\
        );

    \I__1631\ : InMux
    port map (
            O => \N__15639\,
            I => \N__15636\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__15636\,
            I => \N__15633\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__15633\,
            I => \QuadInstance2.un1_Quad_axb_15\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__15630\,
            I => \QuadInstance2.count_enable_cascade_\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__15627\,
            I => \N__15624\
        );

    \I__1626\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15621\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__15621\,
            I => \N__15618\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__15618\,
            I => \QuadInstance2.Quad_RNI1MLE2Z0Z_2\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__15615\,
            I => \QuadInstance2.un1_count_enable_i_a2_0_1_cascade_\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__15612\,
            I => \N__15609\
        );

    \I__1621\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15606\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__15606\,
            I => \N__15603\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__15603\,
            I => \QuadInstance2.Quad_RNI2NLE2Z0Z_3\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__15600\,
            I => \N__15597\
        );

    \I__1617\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15594\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__15594\,
            I => \N__15591\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__15591\,
            I => \QuadInstance2.Quad_RNI4PLE2Z0Z_5\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__15588\,
            I => \N__15585\
        );

    \I__1613\ : InMux
    port map (
            O => \N__15585\,
            I => \N__15582\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__15582\,
            I => \N__15579\
        );

    \I__1611\ : Odrv12
    port map (
            O => \N__15579\,
            I => \QuadInstance2.Quad_RNI5QLE2Z0Z_6\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__15576\,
            I => \N__15571\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__15575\,
            I => \N__15568\
        );

    \I__1608\ : InMux
    port map (
            O => \N__15574\,
            I => \N__15565\
        );

    \I__1607\ : InMux
    port map (
            O => \N__15571\,
            I => \N__15560\
        );

    \I__1606\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15560\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__15565\,
            I => \QuadInstance2.delayedCh_AZ0Z_1\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__15560\,
            I => \QuadInstance2.delayedCh_AZ0Z_1\
        );

    \I__1603\ : InMux
    port map (
            O => \N__15555\,
            I => \N__15552\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__15552\,
            I => \QuadInstance2.delayedCh_AZ0Z_2\
        );

    \I__1601\ : InMux
    port map (
            O => \N__15549\,
            I => \QuadInstance2.un1_Quad_cry_14\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__15546\,
            I => \N__15543\
        );

    \I__1599\ : InMux
    port map (
            O => \N__15543\,
            I => \N__15540\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__15540\,
            I => \QuadInstance2.Quad_RNI8TLE2Z0Z_9\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__15537\,
            I => \N__15534\
        );

    \I__1596\ : InMux
    port map (
            O => \N__15534\,
            I => \N__15531\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__15531\,
            I => \QuadInstance2.Quad_RNIHU2G2Z0Z_11\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \N__15525\
        );

    \I__1593\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15522\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__15522\,
            I => \N__15519\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__15519\,
            I => \QuadInstance2.Quad_RNI0LLE2Z0Z_1\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__15516\,
            I => \N__15513\
        );

    \I__1589\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15510\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__15510\,
            I => \QuadInstance2.Quad_RNIGT2G2Z0Z_10\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__15507\,
            I => \N__15504\
        );

    \I__1586\ : InMux
    port map (
            O => \N__15504\,
            I => \N__15501\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__15501\,
            I => \QuadInstance2.Quad_RNIIV2G2Z0Z_12\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__15498\,
            I => \N__15495\
        );

    \I__1583\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15492\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__15492\,
            I => \N__15489\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__15489\,
            I => \QuadInstance2.Quad_RNI6RLE2Z0Z_7\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__15486\,
            I => \N__15483\
        );

    \I__1579\ : InMux
    port map (
            O => \N__15483\,
            I => \N__15480\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__15480\,
            I => \QuadInstance2.Quad_RNI7SLE2Z0Z_8\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__15477\,
            I => \N__15474\
        );

    \I__1576\ : InMux
    port map (
            O => \N__15474\,
            I => \N__15471\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__15471\,
            I => \N__15468\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__15468\,
            I => \QuadInstance2.Quad_RNI3OLE2Z0Z_4\
        );

    \I__1573\ : InMux
    port map (
            O => \N__15465\,
            I => \QuadInstance2.un1_Quad_cry_5\
        );

    \I__1572\ : InMux
    port map (
            O => \N__15462\,
            I => \QuadInstance2.un1_Quad_cry_6\
        );

    \I__1571\ : InMux
    port map (
            O => \N__15459\,
            I => \bfn_7_7_0_\
        );

    \I__1570\ : InMux
    port map (
            O => \N__15456\,
            I => \QuadInstance2.un1_Quad_cry_8\
        );

    \I__1569\ : InMux
    port map (
            O => \N__15453\,
            I => \QuadInstance2.un1_Quad_cry_9\
        );

    \I__1568\ : InMux
    port map (
            O => \N__15450\,
            I => \QuadInstance2.un1_Quad_cry_10\
        );

    \I__1567\ : InMux
    port map (
            O => \N__15447\,
            I => \QuadInstance2.un1_Quad_cry_11\
        );

    \I__1566\ : InMux
    port map (
            O => \N__15444\,
            I => \QuadInstance2.un1_Quad_cry_12\
        );

    \I__1565\ : InMux
    port map (
            O => \N__15441\,
            I => \QuadInstance2.un1_Quad_cry_13\
        );

    \I__1564\ : InMux
    port map (
            O => \N__15438\,
            I => \N__15435\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__15435\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_15\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__15432\,
            I => \N__15429\
        );

    \I__1561\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15426\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__15426\,
            I => \N__15423\
        );

    \I__1559\ : Span4Mux_h
    port map (
            O => \N__15423\,
            I => \N__15420\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__15420\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_11\
        );

    \I__1557\ : InMux
    port map (
            O => \N__15417\,
            I => \N__15414\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__15414\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_13\
        );

    \I__1555\ : InMux
    port map (
            O => \N__15411\,
            I => \QuadInstance2.un1_Quad_cry_0\
        );

    \I__1554\ : InMux
    port map (
            O => \N__15408\,
            I => \QuadInstance2.un1_Quad_cry_1\
        );

    \I__1553\ : InMux
    port map (
            O => \N__15405\,
            I => \QuadInstance2.un1_Quad_cry_2\
        );

    \I__1552\ : InMux
    port map (
            O => \N__15402\,
            I => \QuadInstance2.un1_Quad_cry_3\
        );

    \I__1551\ : InMux
    port map (
            O => \N__15399\,
            I => \QuadInstance2.un1_Quad_cry_4\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__15396\,
            I => \N__15393\
        );

    \I__1549\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15390\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__15390\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_0\
        );

    \I__1547\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15384\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__15384\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_1\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__15381\,
            I => \N__15378\
        );

    \I__1544\ : InMux
    port map (
            O => \N__15378\,
            I => \N__15375\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__15375\,
            I => \N__15372\
        );

    \I__1542\ : Span4Mux_s3_v
    port map (
            O => \N__15372\,
            I => \N__15369\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__15369\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_7\
        );

    \I__1540\ : InMux
    port map (
            O => \N__15366\,
            I => \N__15363\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__15363\,
            I => \N__15360\
        );

    \I__1538\ : Span4Mux_s3_v
    port map (
            O => \N__15360\,
            I => \N__15357\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__15357\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_8\
        );

    \I__1536\ : InMux
    port map (
            O => \N__15354\,
            I => \N__15351\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__15351\,
            I => \N__15348\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__15348\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_5\
        );

    \I__1533\ : InMux
    port map (
            O => \N__15345\,
            I => \N__15342\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__15342\,
            I => \N__15339\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__15339\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_9\
        );

    \I__1530\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15333\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__15333\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_6\
        );

    \I__1528\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15327\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__15327\,
            I => \N__15324\
        );

    \I__1526\ : Span4Mux_h
    port map (
            O => \N__15324\,
            I => \N__15321\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__15321\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_14\
        );

    \I__1524\ : InMux
    port map (
            O => \N__15318\,
            I => \N__15315\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__15315\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_2\
        );

    \I__1522\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15309\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__15309\,
            I => \N__15306\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__15306\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_3\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__15303\,
            I => \PWMInstance1.un1_periodCounter12_1_0_a2_0_0_cascade_\
        );

    \I__1518\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15297\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__15297\,
            I => \PWMInstance1.PWMPulseWidthCountZ0Z_4\
        );

    \I__1516\ : InMux
    port map (
            O => \N__15294\,
            I => \N__15291\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__15291\,
            I => \N__15288\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__15288\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_1\
        );

    \I__1513\ : InMux
    port map (
            O => \N__15285\,
            I => \N__15282\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__15282\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_0\
        );

    \I__1511\ : CEMux
    port map (
            O => \N__15279\,
            I => \N__15276\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__15276\,
            I => \N__15272\
        );

    \I__1509\ : CEMux
    port map (
            O => \N__15275\,
            I => \N__15267\
        );

    \I__1508\ : Span4Mux_v
    port map (
            O => \N__15272\,
            I => \N__15263\
        );

    \I__1507\ : CEMux
    port map (
            O => \N__15271\,
            I => \N__15260\
        );

    \I__1506\ : CEMux
    port map (
            O => \N__15270\,
            I => \N__15257\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__15267\,
            I => \N__15254\
        );

    \I__1504\ : CEMux
    port map (
            O => \N__15266\,
            I => \N__15251\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__15263\,
            I => \N__15246\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__15260\,
            I => \N__15246\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__15257\,
            I => \N__15243\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__15254\,
            I => \N__15240\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__15251\,
            I => \N__15237\
        );

    \I__1498\ : Span4Mux_v
    port map (
            O => \N__15246\,
            I => \N__15232\
        );

    \I__1497\ : Span4Mux_h
    port map (
            O => \N__15243\,
            I => \N__15232\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__15240\,
            I => \N__15229\
        );

    \I__1495\ : Span4Mux_h
    port map (
            O => \N__15237\,
            I => \N__15226\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__15232\,
            I => \PWMInstance7.pwmWrite_0_7\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__15229\,
            I => \PWMInstance7.pwmWrite_0_7\
        );

    \I__1492\ : Odrv4
    port map (
            O => \N__15226\,
            I => \PWMInstance7.pwmWrite_0_7\
        );

    \I__1491\ : InMux
    port map (
            O => \N__15219\,
            I => \N__15216\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__15216\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_9\
        );

    \I__1489\ : InMux
    port map (
            O => \N__15213\,
            I => \N__15210\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__15210\,
            I => \PWMInstance5.PWMPulseWidthCountZ0Z_8\
        );

    \I__1487\ : IoInMux
    port map (
            O => \N__15207\,
            I => \N__15204\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__15204\,
            I => \RST_c_i\
        );

    \I__1485\ : InMux
    port map (
            O => \N__15201\,
            I => \N__15198\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__15198\,
            I => \ch0_B_c\
        );

    \I__1483\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15192\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__15192\,
            I => \N__15189\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__15189\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_8\
        );

    \I__1480\ : InMux
    port map (
            O => \N__15186\,
            I => \N__15183\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__15183\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_13\
        );

    \I__1478\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15177\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__15177\,
            I => \N__15174\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__15174\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_11\
        );

    \I__1475\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15168\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__15168\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_12\
        );

    \I__1473\ : InMux
    port map (
            O => \N__15165\,
            I => \N__15162\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__15162\,
            I => \N__15159\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__15159\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_5\
        );

    \I__1470\ : InMux
    port map (
            O => \N__15156\,
            I => \N__15153\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__15153\,
            I => \N__15150\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__15150\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_4\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__15147\,
            I => \N__15144\
        );

    \I__1466\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15141\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__15141\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_7\
        );

    \I__1464\ : InMux
    port map (
            O => \N__15138\,
            I => \N__15135\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__15135\,
            I => \N__15132\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__15132\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_6\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__15129\,
            I => \N__15126\
        );

    \I__1460\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15123\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__15123\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_15\
        );

    \I__1458\ : InMux
    port map (
            O => \N__15120\,
            I => \N__15115\
        );

    \I__1457\ : InMux
    port map (
            O => \N__15119\,
            I => \N__15112\
        );

    \I__1456\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15109\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__15115\,
            I => \N__15106\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__15112\,
            I => \N__15103\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__15109\,
            I => \PWMInstance7.periodCounterZ0Z_12\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__15106\,
            I => \PWMInstance7.periodCounterZ0Z_12\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__15103\,
            I => \PWMInstance7.periodCounterZ0Z_12\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__15096\,
            I => \N__15092\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__15095\,
            I => \N__15089\
        );

    \I__1448\ : InMux
    port map (
            O => \N__15092\,
            I => \N__15085\
        );

    \I__1447\ : InMux
    port map (
            O => \N__15089\,
            I => \N__15082\
        );

    \I__1446\ : InMux
    port map (
            O => \N__15088\,
            I => \N__15079\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__15085\,
            I => \N__15074\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__15082\,
            I => \N__15074\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__15079\,
            I => \PWMInstance7.periodCounterZ0Z_13\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__15074\,
            I => \PWMInstance7.periodCounterZ0Z_13\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__15069\,
            I => \N__15066\
        );

    \I__1440\ : InMux
    port map (
            O => \N__15066\,
            I => \N__15063\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__15063\,
            I => \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_6\
        );

    \I__1438\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15057\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__15057\,
            I => \N__15052\
        );

    \I__1436\ : InMux
    port map (
            O => \N__15056\,
            I => \N__15049\
        );

    \I__1435\ : InMux
    port map (
            O => \N__15055\,
            I => \N__15046\
        );

    \I__1434\ : Span4Mux_h
    port map (
            O => \N__15052\,
            I => \N__15043\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__15049\,
            I => \PWMInstance7.periodCounterZ0Z_0\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__15046\,
            I => \PWMInstance7.periodCounterZ0Z_0\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__15043\,
            I => \PWMInstance7.periodCounterZ0Z_0\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__15036\,
            I => \N__15033\
        );

    \I__1429\ : InMux
    port map (
            O => \N__15033\,
            I => \N__15030\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__15030\,
            I => \N__15025\
        );

    \I__1427\ : InMux
    port map (
            O => \N__15029\,
            I => \N__15022\
        );

    \I__1426\ : InMux
    port map (
            O => \N__15028\,
            I => \N__15019\
        );

    \I__1425\ : Span4Mux_h
    port map (
            O => \N__15025\,
            I => \N__15016\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__15022\,
            I => \PWMInstance7.periodCounterZ0Z_1\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__15019\,
            I => \PWMInstance7.periodCounterZ0Z_1\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__15016\,
            I => \PWMInstance7.periodCounterZ0Z_1\
        );

    \I__1421\ : InMux
    port map (
            O => \N__15009\,
            I => \N__15006\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__15006\,
            I => \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_6\
        );

    \I__1419\ : InMux
    port map (
            O => \N__15003\,
            I => \N__15000\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__15000\,
            I => \N__14995\
        );

    \I__1417\ : InMux
    port map (
            O => \N__14999\,
            I => \N__14992\
        );

    \I__1416\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14989\
        );

    \I__1415\ : Span4Mux_h
    port map (
            O => \N__14995\,
            I => \N__14986\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__14992\,
            I => \PWMInstance7.periodCounterZ0Z_6\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__14989\,
            I => \PWMInstance7.periodCounterZ0Z_6\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__14986\,
            I => \PWMInstance7.periodCounterZ0Z_6\
        );

    \I__1411\ : InMux
    port map (
            O => \N__14979\,
            I => \N__14976\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__14976\,
            I => \N__14972\
        );

    \I__1409\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14968\
        );

    \I__1408\ : Span4Mux_h
    port map (
            O => \N__14972\,
            I => \N__14965\
        );

    \I__1407\ : InMux
    port map (
            O => \N__14971\,
            I => \N__14962\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__14968\,
            I => \PWMInstance7.periodCounterZ0Z_7\
        );

    \I__1405\ : Odrv4
    port map (
            O => \N__14965\,
            I => \PWMInstance7.periodCounterZ0Z_7\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__14962\,
            I => \PWMInstance7.periodCounterZ0Z_7\
        );

    \I__1403\ : InMux
    port map (
            O => \N__14955\,
            I => \N__14952\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__14952\,
            I => \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_6\
        );

    \I__1401\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14946\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__14946\,
            I => \N__14943\
        );

    \I__1399\ : Odrv12
    port map (
            O => \N__14943\,
            I => \PWMInstance7.un1_periodCounter12_1_0_a2_0\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__14940\,
            I => \N__14935\
        );

    \I__1397\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14930\
        );

    \I__1396\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14930\
        );

    \I__1395\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14924\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__14930\,
            I => \N__14921\
        );

    \I__1393\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14918\
        );

    \I__1392\ : InMux
    port map (
            O => \N__14928\,
            I => \N__14915\
        );

    \I__1391\ : InMux
    port map (
            O => \N__14927\,
            I => \N__14912\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__14924\,
            I => \N__14909\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__14921\,
            I => \PWMInstance7.out_0_sqmuxa\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__14918\,
            I => \PWMInstance7.out_0_sqmuxa\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__14915\,
            I => \PWMInstance7.out_0_sqmuxa\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__14912\,
            I => \PWMInstance7.out_0_sqmuxa\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__14909\,
            I => \PWMInstance7.out_0_sqmuxa\
        );

    \I__1384\ : InMux
    port map (
            O => \N__14898\,
            I => \bfn_3_11_0_\
        );

    \I__1383\ : IoInMux
    port map (
            O => \N__14895\,
            I => \N__14892\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__14892\,
            I => \N__14889\
        );

    \I__1381\ : Span4Mux_s3_v
    port map (
            O => \N__14889\,
            I => \N__14886\
        );

    \I__1380\ : Span4Mux_h
    port map (
            O => \N__14886\,
            I => \N__14883\
        );

    \I__1379\ : Span4Mux_v
    port map (
            O => \N__14883\,
            I => \N__14879\
        );

    \I__1378\ : InMux
    port map (
            O => \N__14882\,
            I => \N__14876\
        );

    \I__1377\ : Odrv4
    port map (
            O => \N__14879\,
            I => \PWM7_c\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__14876\,
            I => \PWM7_c\
        );

    \I__1375\ : InMux
    port map (
            O => \N__14871\,
            I => \N__14865\
        );

    \I__1374\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14865\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__14865\,
            I => \pwmWrite_fastZ0Z_7\
        );

    \I__1372\ : InMux
    port map (
            O => \N__14862\,
            I => \N__14859\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__14859\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_9\
        );

    \I__1370\ : InMux
    port map (
            O => \N__14856\,
            I => \N__14853\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__14853\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_10\
        );

    \I__1368\ : InMux
    port map (
            O => \N__14850\,
            I => \N__14847\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__14847\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_3\
        );

    \I__1366\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14839\
        );

    \I__1365\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14836\
        );

    \I__1364\ : InMux
    port map (
            O => \N__14842\,
            I => \N__14833\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__14839\,
            I => \N__14828\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__14836\,
            I => \N__14828\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__14833\,
            I => \N__14825\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__14828\,
            I => \PWMInstance7.periodCounterZ0Z_15\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__14825\,
            I => \PWMInstance7.periodCounterZ0Z_15\
        );

    \I__1358\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14816\
        );

    \I__1357\ : InMux
    port map (
            O => \N__14819\,
            I => \N__14813\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__14816\,
            I => \N__14807\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__14813\,
            I => \N__14807\
        );

    \I__1354\ : InMux
    port map (
            O => \N__14812\,
            I => \N__14804\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__14807\,
            I => \PWMInstance7.periodCounterZ0Z_14\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__14804\,
            I => \PWMInstance7.periodCounterZ0Z_14\
        );

    \I__1351\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14796\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__14796\,
            I => \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_6\
        );

    \I__1349\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14790\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__14790\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_14\
        );

    \I__1347\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14782\
        );

    \I__1346\ : InMux
    port map (
            O => \N__14786\,
            I => \N__14777\
        );

    \I__1345\ : InMux
    port map (
            O => \N__14785\,
            I => \N__14777\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__14782\,
            I => \PWMInstance7.periodCounterZ0Z_4\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__14777\,
            I => \PWMInstance7.periodCounterZ0Z_4\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__14772\,
            I => \N__14767\
        );

    \I__1341\ : InMux
    port map (
            O => \N__14771\,
            I => \N__14764\
        );

    \I__1340\ : InMux
    port map (
            O => \N__14770\,
            I => \N__14759\
        );

    \I__1339\ : InMux
    port map (
            O => \N__14767\,
            I => \N__14759\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__14764\,
            I => \PWMInstance7.periodCounterZ0Z_5\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__14759\,
            I => \PWMInstance7.periodCounterZ0Z_5\
        );

    \I__1336\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14749\
        );

    \I__1335\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14744\
        );

    \I__1334\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14744\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__14749\,
            I => \PWMInstance7.periodCounterZ0Z_8\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__14744\,
            I => \PWMInstance7.periodCounterZ0Z_8\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__14739\,
            I => \N__14734\
        );

    \I__1330\ : InMux
    port map (
            O => \N__14738\,
            I => \N__14731\
        );

    \I__1329\ : InMux
    port map (
            O => \N__14737\,
            I => \N__14726\
        );

    \I__1328\ : InMux
    port map (
            O => \N__14734\,
            I => \N__14726\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__14731\,
            I => \PWMInstance7.periodCounterZ0Z_9\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__14726\,
            I => \PWMInstance7.periodCounterZ0Z_9\
        );

    \I__1325\ : InMux
    port map (
            O => \N__14721\,
            I => \N__14718\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__14718\,
            I => \N__14715\
        );

    \I__1323\ : Odrv12
    port map (
            O => \N__14715\,
            I => \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_6\
        );

    \I__1322\ : InMux
    port map (
            O => \N__14712\,
            I => \N__14709\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__14709\,
            I => \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_6\
        );

    \I__1320\ : InMux
    port map (
            O => \N__14706\,
            I => \N__14703\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__14703\,
            I => \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_6\
        );

    \I__1318\ : InMux
    port map (
            O => \N__14700\,
            I => \N__14697\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__14697\,
            I => \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_6\
        );

    \I__1316\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14682\
        );

    \I__1315\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14682\
        );

    \I__1314\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14682\
        );

    \I__1313\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14682\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__14682\,
            I => \PWMInstance7.clkCountZ0Z_0\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__14679\,
            I => \N__14675\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__14678\,
            I => \N__14672\
        );

    \I__1309\ : InMux
    port map (
            O => \N__14675\,
            I => \N__14661\
        );

    \I__1308\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14661\
        );

    \I__1307\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14661\
        );

    \I__1306\ : InMux
    port map (
            O => \N__14670\,
            I => \N__14661\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__14661\,
            I => \PWMInstance7.clkCountZ0Z_1\
        );

    \I__1304\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14655\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__14655\,
            I => \PWMInstance7.PWMPulseWidthCountZ0Z_2\
        );

    \I__1302\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14647\
        );

    \I__1301\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14642\
        );

    \I__1300\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14642\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__14647\,
            I => \PWMInstance7.periodCounterZ0Z_2\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__14642\,
            I => \PWMInstance7.periodCounterZ0Z_2\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__14637\,
            I => \N__14632\
        );

    \I__1296\ : InMux
    port map (
            O => \N__14636\,
            I => \N__14629\
        );

    \I__1295\ : InMux
    port map (
            O => \N__14635\,
            I => \N__14626\
        );

    \I__1294\ : InMux
    port map (
            O => \N__14632\,
            I => \N__14623\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__14629\,
            I => \PWMInstance7.periodCounterZ0Z_3\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__14626\,
            I => \PWMInstance7.periodCounterZ0Z_3\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__14623\,
            I => \PWMInstance7.periodCounterZ0Z_3\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__14616\,
            I => \N__14612\
        );

    \I__1289\ : InMux
    port map (
            O => \N__14615\,
            I => \N__14608\
        );

    \I__1288\ : InMux
    port map (
            O => \N__14612\,
            I => \N__14603\
        );

    \I__1287\ : InMux
    port map (
            O => \N__14611\,
            I => \N__14603\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__14608\,
            I => \PWMInstance7.periodCounterZ0Z_11\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__14603\,
            I => \PWMInstance7.periodCounterZ0Z_11\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__14598\,
            I => \N__14593\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__14597\,
            I => \N__14590\
        );

    \I__1282\ : InMux
    port map (
            O => \N__14596\,
            I => \N__14587\
        );

    \I__1281\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14582\
        );

    \I__1280\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14582\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__14587\,
            I => \PWMInstance7.periodCounterZ0Z_10\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__14582\,
            I => \PWMInstance7.periodCounterZ0Z_10\
        );

    \I__1277\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14574\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__14574\,
            I => \PWMInstance7.un1_periodCounter12_1_0_a2_0_0\
        );

    \I__1275\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14568\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__14568\,
            I => \PWMInstance7.un1_periodCounter12_1_0_a2_0_10\
        );

    \I__1273\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14562\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__14562\,
            I => \PWMInstance7.un1_periodCounter12_1_0_a2_0_9\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__14559\,
            I => \PWMInstance7.un1_periodCounter12_1_0_a2_0_12_cascade_\
        );

    \I__1270\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14553\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__14553\,
            I => \N__14550\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__14550\,
            I => \PWMInstance7.un1_periodCounter12_1_0_a2_0_14\
        );

    \I__1267\ : InMux
    port map (
            O => \N__14547\,
            I => \PWMInstance7.un1_periodCounter_2_cry_10\
        );

    \I__1266\ : InMux
    port map (
            O => \N__14544\,
            I => \PWMInstance7.un1_periodCounter_2_cry_11\
        );

    \I__1265\ : InMux
    port map (
            O => \N__14541\,
            I => \PWMInstance7.un1_periodCounter_2_cry_12\
        );

    \I__1264\ : InMux
    port map (
            O => \N__14538\,
            I => \PWMInstance7.un1_periodCounter_2_cry_13\
        );

    \I__1263\ : InMux
    port map (
            O => \N__14535\,
            I => \PWMInstance7.un1_periodCounter_2_cry_14\
        );

    \I__1262\ : InMux
    port map (
            O => \N__14532\,
            I => \bfn_2_10_0_\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__14529\,
            I => \N__14526\
        );

    \I__1260\ : InMux
    port map (
            O => \N__14526\,
            I => \N__14521\
        );

    \I__1259\ : InMux
    port map (
            O => \N__14525\,
            I => \N__14518\
        );

    \I__1258\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14515\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__14521\,
            I => \N__14512\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__14518\,
            I => \N__14509\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__14515\,
            I => \PWMInstance7.periodCounterZ0Z_16\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__14512\,
            I => \PWMInstance7.periodCounterZ0Z_16\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__14509\,
            I => \PWMInstance7.periodCounterZ0Z_16\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__14502\,
            I => \N__14498\
        );

    \I__1251\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14494\
        );

    \I__1250\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14491\
        );

    \I__1249\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14488\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__14494\,
            I => \PWMInstance7.periodCounter12\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__14491\,
            I => \PWMInstance7.periodCounter12\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__14488\,
            I => \PWMInstance7.periodCounter12\
        );

    \I__1245\ : InMux
    port map (
            O => \N__14481\,
            I => \PWMInstance7.un1_periodCounter_2_cry_1\
        );

    \I__1244\ : InMux
    port map (
            O => \N__14478\,
            I => \PWMInstance7.un1_periodCounter_2_cry_2\
        );

    \I__1243\ : InMux
    port map (
            O => \N__14475\,
            I => \PWMInstance7.un1_periodCounter_2_cry_3\
        );

    \I__1242\ : InMux
    port map (
            O => \N__14472\,
            I => \PWMInstance7.un1_periodCounter_2_cry_4\
        );

    \I__1241\ : InMux
    port map (
            O => \N__14469\,
            I => \PWMInstance7.un1_periodCounter_2_cry_5\
        );

    \I__1240\ : InMux
    port map (
            O => \N__14466\,
            I => \PWMInstance7.un1_periodCounter_2_cry_6\
        );

    \I__1239\ : InMux
    port map (
            O => \N__14463\,
            I => \bfn_2_9_0_\
        );

    \I__1238\ : InMux
    port map (
            O => \N__14460\,
            I => \PWMInstance7.un1_periodCounter_2_cry_8\
        );

    \I__1237\ : InMux
    port map (
            O => \N__14457\,
            I => \PWMInstance7.un1_periodCounter_2_cry_9\
        );

    \I__1236\ : IoInMux
    port map (
            O => \N__14454\,
            I => \N__14451\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__14451\,
            I => \N__14448\
        );

    \I__1234\ : IoSpan4Mux
    port map (
            O => \N__14448\,
            I => \N__14445\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__14445\,
            I => \CLK_c\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__14442\,
            I => \PWMInstance7.un1_periodCounter12_1_0_a2_0_6_cascade_\
        );

    \I__1231\ : InMux
    port map (
            O => \N__14439\,
            I => \PWMInstance7.un1_periodCounter_2_cry_0\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \QuadInstance7.un1_Quad_cry_7\,
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \QuadInstance6.un1_Quad_cry_7\,
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_10_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_6_0_\
        );

    \IN_MUX_bfv_10_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \QuadInstance5.un1_Quad_cry_7\,
            carryinitout => \bfn_10_7_0_\
        );

    \IN_MUX_bfv_15_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_3_0_\
        );

    \IN_MUX_bfv_15_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \QuadInstance4.un1_Quad_cry_7\,
            carryinitout => \bfn_15_4_0_\
        );

    \IN_MUX_bfv_10_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_8_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \QuadInstance3.un1_Quad_cry_7\,
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \QuadInstance2.un1_Quad_cry_7\,
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \QuadInstance1.un1_Quad_cry_7\,
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_17_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_6_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \QuadInstance0.un1_Quad_cry_7\,
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_3_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_10_0_\
        );

    \IN_MUX_bfv_3_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_7\,
            carryinitout => \bfn_3_11_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_7\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_7\,
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_15_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_1_0_\
        );

    \IN_MUX_bfv_15_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_7\,
            carryinitout => \bfn_15_2_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_7\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_7\,
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_7\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_7\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance7.un1_periodCounter_2_cry_7\,
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance7.un1_periodCounter_2_cry_15\,
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance6.un1_periodCounter_2_cry_7\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance6.un1_periodCounter_2_cry_15\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance5.un1_periodCounter_2_cry_7\,
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance5.un1_periodCounter_2_cry_15\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance4.un1_periodCounter_2_cry_7\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance4.un1_periodCounter_2_cry_15\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance3.un1_periodCounter_2_cry_7\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance3.un1_periodCounter_2_cry_15\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance2.un1_periodCounter_2_cry_7\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance2.un1_periodCounter_2_cry_15\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance1.un1_periodCounter_2_cry_7\,
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance1.un1_periodCounter_2_cry_15\,
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance0.un1_periodCounter_2_cry_7\,
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_7_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWMInstance0.un1_periodCounter_2_cry_15\,
            carryinitout => \bfn_7_18_0_\
        );

    \internalOscilator\ : SMCCLK
    port map (
            CLK => \internalOscilatorOutputNet\
        );

    \SCKr_RNIBA7C_0_2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__37941\,
            GLOBALBUFFEROUTPUT => \N_1187_g\
        );

    \SCKr_RNIMKEO_0_2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__37923\,
            GLOBALBUFFEROUTPUT => \N_45_0_g\
        );

    \RST_ibuf_RNIUR47_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__15207\,
            GLOBALBUFFEROUTPUT => \RST_c_i_g\
        );

    \PWMInstance0.N_42_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__25626\,
            GLOBALBUFFEROUTPUT => \PWMInstance0_N_42_g\
        );

    \My_Global_Buffer_i\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14454\,
            GLOBALBUFFEROUTPUT => myclk
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PWMInstance7.periodCounter_RNIG0CG_16_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14525\,
            in2 => \_gnd_net_\,
            in3 => \N__14971\,
            lcout => OPEN,
            ltout => \PWMInstance7.un1_periodCounter12_1_0_a2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.periodCounter_RNI7VP12_1_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14842\,
            in1 => \N__15028\,
            in2 => \N__14442\,
            in3 => \N__14497\,
            lcout => \PWMInstance7.un1_periodCounter12_1_0_a2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.periodCounter_0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15055\,
            in2 => \N__14502\,
            in3 => \N__14501\,
            lcout => \PWMInstance7.periodCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_0\,
            clk => \N__38625\,
            ce => 'H',
            sr => \N__35314\
        );

    \PWMInstance7.periodCounter_1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15029\,
            in2 => \_gnd_net_\,
            in3 => \N__14439\,
            lcout => \PWMInstance7.periodCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_0\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_1\,
            clk => \N__38625\,
            ce => 'H',
            sr => \N__35314\
        );

    \PWMInstance7.periodCounter_2_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14652\,
            in2 => \_gnd_net_\,
            in3 => \N__14481\,
            lcout => \PWMInstance7.periodCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_1\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_2\,
            clk => \N__38625\,
            ce => 'H',
            sr => \N__35314\
        );

    \PWMInstance7.periodCounter_3_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14636\,
            in2 => \_gnd_net_\,
            in3 => \N__14478\,
            lcout => \PWMInstance7.periodCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_2\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_3\,
            clk => \N__38625\,
            ce => 'H',
            sr => \N__35314\
        );

    \PWMInstance7.periodCounter_4_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14787\,
            in2 => \_gnd_net_\,
            in3 => \N__14475\,
            lcout => \PWMInstance7.periodCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_3\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_4\,
            clk => \N__38625\,
            ce => 'H',
            sr => \N__35314\
        );

    \PWMInstance7.periodCounter_5_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14771\,
            in2 => \_gnd_net_\,
            in3 => \N__14472\,
            lcout => \PWMInstance7.periodCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_4\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_5\,
            clk => \N__38625\,
            ce => 'H',
            sr => \N__35314\
        );

    \PWMInstance7.periodCounter_6_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14999\,
            in2 => \_gnd_net_\,
            in3 => \N__14469\,
            lcout => \PWMInstance7.periodCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_5\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_6\,
            clk => \N__38625\,
            ce => 'H',
            sr => \N__35314\
        );

    \PWMInstance7.periodCounter_7_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14929\,
            in1 => \N__14975\,
            in2 => \_gnd_net_\,
            in3 => \N__14466\,
            lcout => \PWMInstance7.periodCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_6\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_7\,
            clk => \N__38625\,
            ce => 'H',
            sr => \N__35314\
        );

    \PWMInstance7.periodCounter_8_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14754\,
            in2 => \_gnd_net_\,
            in3 => \N__14463\,
            lcout => \PWMInstance7.periodCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_8\,
            clk => \N__38614\,
            ce => 'H',
            sr => \N__35312\
        );

    \PWMInstance7.periodCounter_9_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14738\,
            in2 => \_gnd_net_\,
            in3 => \N__14460\,
            lcout => \PWMInstance7.periodCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_8\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_9\,
            clk => \N__38614\,
            ce => 'H',
            sr => \N__35312\
        );

    \PWMInstance7.periodCounter_10_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14596\,
            in2 => \_gnd_net_\,
            in3 => \N__14457\,
            lcout => \PWMInstance7.periodCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_9\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_10\,
            clk => \N__38614\,
            ce => 'H',
            sr => \N__35312\
        );

    \PWMInstance7.periodCounter_11_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14938\,
            in1 => \N__14615\,
            in2 => \_gnd_net_\,
            in3 => \N__14547\,
            lcout => \PWMInstance7.periodCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_10\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_11\,
            clk => \N__38614\,
            ce => 'H',
            sr => \N__35312\
        );

    \PWMInstance7.periodCounter_12_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14927\,
            in1 => \N__15118\,
            in2 => \_gnd_net_\,
            in3 => \N__14544\,
            lcout => \PWMInstance7.periodCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_11\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_12\,
            clk => \N__38614\,
            ce => 'H',
            sr => \N__35312\
        );

    \PWMInstance7.periodCounter_13_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14939\,
            in1 => \N__15088\,
            in2 => \_gnd_net_\,
            in3 => \N__14541\,
            lcout => \PWMInstance7.periodCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_12\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_13\,
            clk => \N__38614\,
            ce => 'H',
            sr => \N__35312\
        );

    \PWMInstance7.periodCounter_14_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14820\,
            in2 => \_gnd_net_\,
            in3 => \N__14538\,
            lcout => \PWMInstance7.periodCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_13\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_14\,
            clk => \N__38614\,
            ce => 'H',
            sr => \N__35312\
        );

    \PWMInstance7.periodCounter_15_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14844\,
            in2 => \_gnd_net_\,
            in3 => \N__14535\,
            lcout => \PWMInstance7.periodCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_periodCounter_2_cry_14\,
            carryout => \PWMInstance7.un1_periodCounter_2_cry_15\,
            clk => \N__38614\,
            ce => 'H',
            sr => \N__35312\
        );

    \PWMInstance7.periodCounter_16_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14928\,
            in1 => \N__14524\,
            in2 => \_gnd_net_\,
            in3 => \N__14532\,
            lcout => \PWMInstance7.periodCounterZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38603\,
            ce => 'H',
            sr => \N__35311\
        );

    \PWMInstance7.out_RNO_0_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__14871\,
            in1 => \N__14671\,
            in2 => \N__14529\,
            in3 => \N__14692\,
            lcout => \PWMInstance7.un1_periodCounter12_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.clkCount_0_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000101"
        )
    port map (
            in0 => \N__14693\,
            in1 => \_gnd_net_\,
            in2 => \N__14678\,
            in3 => \N__17813\,
            lcout => \PWMInstance7.clkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38626\,
            ce => 'H',
            sr => \N__35695\
        );

    \PWMInstance7.clkCount_RNIE5211_0_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__14870\,
            in1 => \N__14670\,
            in2 => \_gnd_net_\,
            in3 => \N__14691\,
            lcout => \PWMInstance7.periodCounter12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.clkCount_1_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000001010"
        )
    port map (
            in0 => \N__14694\,
            in1 => \_gnd_net_\,
            in2 => \N__14679\,
            in3 => \N__17814\,
            lcout => \PWMInstance7.clkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38626\,
            ce => 'H',
            sr => \N__35695\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__14651\,
            in1 => \N__14850\,
            in2 => \N__14637\,
            in3 => \N__14658\,
            lcout => \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_2_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31604\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38615\,
            ce => \N__15270\,
            sr => \N__35702\
        );

    \PWMInstance7.periodCounter_RNI9PBG_2_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14812\,
            in2 => \_gnd_net_\,
            in3 => \N__14650\,
            lcout => \PWMInstance7.un1_periodCounter12_1_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.periodCounter_RNI79MR_3_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14737\,
            in1 => \N__14770\,
            in2 => \N__14616\,
            in3 => \N__14635\,
            lcout => \PWMInstance7.un1_periodCounter12_1_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__15180\,
            in1 => \N__14611\,
            in2 => \N__14597\,
            in3 => \N__14856\,
            lcout => \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.periodCounter_RNI68MR_0_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14753\,
            in1 => \N__14998\,
            in2 => \N__15095\,
            in3 => \N__15056\,
            lcout => \PWMInstance7.un1_periodCounter12_1_0_a2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.periodCounter_RNIS3EB1_4_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14786\,
            in1 => \N__15120\,
            in2 => \N__14598\,
            in3 => \N__14577\,
            lcout => OPEN,
            ltout => \PWMInstance7.un1_periodCounter12_1_0_a2_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.periodCounter_RNIGKK45_0_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14571\,
            in1 => \N__14565\,
            in2 => \N__14559\,
            in3 => \N__14556\,
            lcout => \PWMInstance7.out_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__14785\,
            in1 => \N__15165\,
            in2 => \N__14772\,
            in3 => \N__15156\,
            lcout => \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__14752\,
            in1 => \N__14862\,
            in2 => \N__14739\,
            in3 => \N__15195\,
            lcout => \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15009\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_10_0_\,
            carryout => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14721\,
            in2 => \N__32585\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_0\,
            carryout => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14712\,
            in2 => \N__32580\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_1\,
            carryout => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14955\,
            in2 => \N__32583\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_2\,
            carryout => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14706\,
            in2 => \N__32581\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_3\,
            carryout => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14700\,
            in2 => \N__32584\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_4\,
            carryout => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32534\,
            in2 => \N__15069\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_5\,
            carryout => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14799\,
            in2 => \N__32582\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_6\,
            carryout => \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.out_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__14882\,
            in1 => \N__14949\,
            in2 => \N__14940\,
            in3 => \N__14898\,
            lcout => \PWM7_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38585\,
            ce => 'H',
            sr => \N__35726\
        );

    \pwmWrite_fast_7_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__33857\,
            in1 => \N__33670\,
            in2 => \N__33449\,
            in3 => \N__23463\,
            lcout => \pwmWrite_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_9_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28580\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38604\,
            ce => \N__15266\,
            sr => \N__35696\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_10_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36167\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38604\,
            ce => \N__15266\,
            sr => \N__35696\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_3_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32084\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38604\,
            ce => \N__15266\,
            sr => \N__35696\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__14793\,
            in1 => \N__14843\,
            in2 => \N__15129\,
            in3 => \N__14819\,
            lcout => \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_14_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34399\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38595\,
            ce => \N__15279\,
            sr => \N__35703\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__15171\,
            in1 => \N__15119\,
            in2 => \N__15096\,
            in3 => \N__15186\,
            lcout => \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__15294\,
            in1 => \N__15060\,
            in2 => \N__15036\,
            in3 => \N__15285\,
            lcout => \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__15003\,
            in1 => \N__15138\,
            in2 => \N__15147\,
            in3 => \N__14979\,
            lcout => \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_10_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36166\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38557\,
            ce => \N__19651\,
            sr => \N__35736\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_9_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28579\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38551\,
            ce => \N__19653\,
            sr => \N__35741\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_8_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29007\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38637\,
            ce => \N__16826\,
            sr => \N__35678\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_7_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29417\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38637\,
            ce => \N__16826\,
            sr => \N__35678\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_11_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36003\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38637\,
            ce => \N__16826\,
            sr => \N__35678\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_14_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34414\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38605\,
            ce => \N__16822\,
            sr => \N__35683\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_ctle_15_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__35824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17807\,
            lcout => \PWMInstance7.pwmWrite_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_8_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29003\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38586\,
            ce => \N__15275\,
            sr => \N__35697\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_13_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28725\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38586\,
            ce => \N__15275\,
            sr => \N__35697\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_11_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36002\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38586\,
            ce => \N__15275\,
            sr => \N__35697\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_12_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28873\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38586\,
            ce => \N__15275\,
            sr => \N__35697\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_5_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36376\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38586\,
            ce => \N__15275\,
            sr => \N__35697\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_4_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36503\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38586\,
            ce => \N__15275\,
            sr => \N__35697\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_7_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29460\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38574\,
            ce => \N__15271\,
            sr => \N__35704\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_6_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31125\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38574\,
            ce => \N__15271\,
            sr => \N__35704\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_15_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31894\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38574\,
            ce => \N__15271\,
            sr => \N__35704\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_1_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31278\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38574\,
            ce => \N__15271\,
            sr => \N__35704\
        );

    \PWMInstance7.PWMPulseWidthCount_esr_0_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31436\,
            lcout => \PWMInstance7.PWMPulseWidthCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38574\,
            ce => \N__15271\,
            sr => \N__35704\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_10_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36149\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38565\,
            ce => \N__18249\,
            sr => \N__35708\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_8_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29002\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38558\,
            ce => \N__19650\,
            sr => \N__35718\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_14_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34413\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38558\,
            ce => \N__19650\,
            sr => \N__35718\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__17942\,
            in1 => \N__15219\,
            in2 => \N__19419\,
            in3 => \N__15213\,
            lcout => \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_12_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28872\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38547\,
            ce => \N__19652\,
            sr => \N__35737\
        );

    \RST_ibuf_RNIUR47_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34515\,
            lcout => \RST_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.delayedCh_B_0_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15201\,
            lcout => \QuadInstance0.delayedCh_BZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.periodCounter_RNIFA3I1_3_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16201\,
            in1 => \N__16129\,
            in2 => \N__16349\,
            in3 => \N__16240\,
            lcout => \PWMInstance1.un1_periodCounter12_1_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__16022\,
            in1 => \N__15312\,
            in2 => \N__16242\,
            in3 => \N__15318\,
            lcout => \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_2_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31608\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38658\,
            ce => \N__16827\,
            sr => \N__35676\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_3_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32091\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38658\,
            ce => \N__16827\,
            sr => \N__35676\
        );

    \PWMInstance1.periodCounter_RNIT6VP_2_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16267\,
            in2 => \_gnd_net_\,
            in3 => \N__16021\,
            lcout => OPEN,
            ltout => \PWMInstance1.un1_periodCounter12_1_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.periodCounter_RNIUIR12_4_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16318\,
            in1 => \N__16102\,
            in2 => \N__15303\,
            in3 => \N__16220\,
            lcout => \PWMInstance1.un1_periodCounter12_1_0_a2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__16219\,
            in1 => \N__15354\,
            in2 => \N__16203\,
            in3 => \N__15300\,
            lcout => \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_4_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38658\,
            ce => \N__16827\,
            sr => \N__35676\
        );

    \PWMInstance1.periodCounter_RNIE93I1_0_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16044\,
            in1 => \N__16295\,
            in2 => \N__16182\,
            in3 => \N__16151\,
            lcout => \PWMInstance1.un1_periodCounter12_1_0_a2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__15387\,
            in1 => \N__16043\,
            in2 => \N__15396\,
            in3 => \N__16619\,
            lcout => \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_0_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31435\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38648\,
            ce => \N__16823\,
            sr => \N__35677\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_1_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31279\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38648\,
            ce => \N__16823\,
            sr => \N__35677\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__16178\,
            in1 => \N__15336\,
            in2 => \N__15381\,
            in3 => \N__16682\,
            lcout => \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__15345\,
            in1 => \N__16150\,
            in2 => \N__16131\,
            in3 => \N__15366\,
            lcout => \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_13_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28728\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38638\,
            ce => \N__16825\,
            sr => \N__35679\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_5_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36377\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38638\,
            ce => \N__16825\,
            sr => \N__35679\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_9_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28584\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38638\,
            ce => \N__16825\,
            sr => \N__35679\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_6_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31124\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38638\,
            ce => \N__16825\,
            sr => \N__35679\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__15438\,
            in1 => \N__15330\,
            in2 => \N__16659\,
            in3 => \N__16272\,
            lcout => \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_15_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31918\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38627\,
            ce => \N__16824\,
            sr => \N__35680\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__16107\,
            in1 => \N__16365\,
            in2 => \N__15432\,
            in3 => \N__16350\,
            lcout => \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__16323\,
            in1 => \N__16299\,
            in2 => \N__16374\,
            in3 => \N__15417\,
            lcout => \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.un1_Quad_cry_0_c_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18529\,
            in2 => \N__30845\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \QuadInstance2.un1_Quad_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23834\,
            in2 => \N__15528\,
            in3 => \N__15411\,
            lcout => \QuadInstance2.Quad_RNO_0_1_1\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_0\,
            carryout => \QuadInstance2.un1_Quad_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30461\,
            in2 => \N__15627\,
            in3 => \N__15408\,
            lcout => \QuadInstance2.Quad_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_1\,
            carryout => \QuadInstance2.un1_Quad_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24406\,
            in2 => \N__15612\,
            in3 => \N__15405\,
            lcout => \QuadInstance2.Quad_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_2\,
            carryout => \QuadInstance2.un1_Quad_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_4_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21296\,
            in2 => \N__15477\,
            in3 => \N__15402\,
            lcout => \QuadInstance2.Quad_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_3\,
            carryout => \QuadInstance2.un1_Quad_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_5_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23717\,
            in2 => \N__15600\,
            in3 => \N__15399\,
            lcout => \QuadInstance2.Quad_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_4\,
            carryout => \QuadInstance2.un1_Quad_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_6_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28300\,
            in2 => \N__15588\,
            in3 => \N__15465\,
            lcout => \QuadInstance2.Quad_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_5\,
            carryout => \QuadInstance2.un1_Quad_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_7_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26374\,
            in2 => \N__15498\,
            in3 => \N__15462\,
            lcout => \QuadInstance2.Quad_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_6\,
            carryout => \QuadInstance2.un1_Quad_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_8_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30703\,
            in2 => \N__15486\,
            in3 => \N__15459\,
            lcout => \QuadInstance2.Quad_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \QuadInstance2.un1_Quad_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_9_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25438\,
            in2 => \N__15546\,
            in3 => \N__15456\,
            lcout => \QuadInstance2.Quad_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_8\,
            carryout => \QuadInstance2.un1_Quad_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_10_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34675\,
            in2 => \N__15516\,
            in3 => \N__15453\,
            lcout => \QuadInstance2.Quad_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_9\,
            carryout => \QuadInstance2.un1_Quad_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_11_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22451\,
            in2 => \N__15537\,
            in3 => \N__15450\,
            lcout => \QuadInstance2.Quad_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_10\,
            carryout => \QuadInstance2.un1_Quad_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_12_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22351\,
            in2 => \N__15507\,
            in3 => \N__15447\,
            lcout => \QuadInstance2.Quad_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_11\,
            carryout => \QuadInstance2.un1_Quad_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_13_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19973\,
            in2 => \N__17520\,
            in3 => \N__15444\,
            lcout => \QuadInstance2.Quad_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_12\,
            carryout => \QuadInstance2.un1_Quad_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_14_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15714\,
            in2 => \N__20047\,
            in3 => \N__15441\,
            lcout => \QuadInstance2.Quad_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \QuadInstance2.un1_Quad_cry_13\,
            carryout => \QuadInstance2.un1_Quad_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_15_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__15639\,
            in1 => \N__22159\,
            in2 => \N__31923\,
            in3 => \N__15549\,
            lcout => \dataRead2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38606\,
            ce => 'H',
            sr => \N__35684\
        );

    \QuadInstance2.Quad_RNI8TLE2_9_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__25442\,
            in1 => \N__22102\,
            in2 => \N__18518\,
            in3 => \N__17572\,
            lcout => \QuadInstance2.Quad_RNI8TLE2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNIHU2G2_11_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__22105\,
            in1 => \N__22455\,
            in2 => \N__17592\,
            in3 => \N__18503\,
            lcout => \QuadInstance2.Quad_RNIHU2G2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNI0LLE2_1_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__23835\,
            in1 => \N__22098\,
            in2 => \N__18516\,
            in3 => \N__17561\,
            lcout => \QuadInstance2.Quad_RNI0LLE2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNIGT2G2_10_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__22103\,
            in1 => \N__34676\,
            in2 => \N__17591\,
            in3 => \N__18499\,
            lcout => \QuadInstance2.Quad_RNIGT2G2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNIIV2G2_12_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__22352\,
            in1 => \N__22104\,
            in2 => \N__18519\,
            in3 => \N__17576\,
            lcout => \QuadInstance2.Quad_RNIIV2G2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNI6RLE2_7_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__22100\,
            in1 => \N__26375\,
            in2 => \N__17590\,
            in3 => \N__18492\,
            lcout => \QuadInstance2.Quad_RNI6RLE2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNI7SLE2_8_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__30711\,
            in1 => \N__22101\,
            in2 => \N__18517\,
            in3 => \N__17568\,
            lcout => \QuadInstance2.Quad_RNI7SLE2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNI3OLE2_4_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__22099\,
            in1 => \N__21297\,
            in2 => \N__17589\,
            in3 => \N__18491\,
            lcout => \QuadInstance2.Quad_RNI3OLE2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNO_0_15_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111110000"
        )
    port map (
            in0 => \N__22110\,
            in1 => \N__17584\,
            in2 => \N__24314\,
            in3 => \N__18507\,
            lcout => \QuadInstance2.un1_Quad_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.delayedCh_A_RNIK9UB1_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15555\,
            in1 => \N__15693\,
            in2 => \N__15575\,
            in3 => \N__15704\,
            lcout => \QuadInstance2.count_enable\,
            ltout => \QuadInstance2.count_enable_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNI1MLE2_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__22106\,
            in1 => \N__30465\,
            in2 => \N__15630\,
            in3 => \N__17577\,
            lcout => \QuadInstance2.Quad_RNI1MLE2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.delayedCh_B_RNIO04T_2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__34471\,
            in1 => \_gnd_net_\,
            in2 => \N__15576\,
            in3 => \N__15692\,
            lcout => \QuadInstance2.un1_count_enable_i_a2_0_1\,
            ltout => \QuadInstance2.un1_count_enable_i_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNI2NLE2_3_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__22107\,
            in1 => \N__24414\,
            in2 => \N__15615\,
            in3 => \N__18504\,
            lcout => \QuadInstance2.Quad_RNI2NLE2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNI4PLE2_5_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001010"
        )
    port map (
            in0 => \N__18506\,
            in1 => \N__22109\,
            in2 => \N__17594\,
            in3 => \N__23718\,
            lcout => \QuadInstance2.Quad_RNI4PLE2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_15_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111001100"
        )
    port map (
            in0 => \N__16522\,
            in1 => \N__24290\,
            in2 => \N__26011\,
            in3 => \N__21795\,
            lcout => \QuadInstance7.un1_Quad_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNI5QLE2_6_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001010"
        )
    port map (
            in0 => \N__18505\,
            in1 => \N__22108\,
            in2 => \N__17593\,
            in3 => \N__28305\,
            lcout => \QuadInstance2.Quad_RNI5QLE2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.delayedCh_A_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance2.delayedCh_AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.delayedCh_A_2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15574\,
            lcout => \QuadInstance2.delayedCh_AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.delayedCh_B_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23313\,
            lcout => \QuadInstance2.delayedCh_BZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNIK13G2_14_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__22150\,
            in1 => \N__18515\,
            in2 => \N__20049\,
            in3 => \N__17588\,
            lcout => \QuadInstance2.Quad_RNIK13G2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.delayedCh_B_2_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15705\,
            lcout => \QuadInstance2.delayedCh_BZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_fast_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__33846\,
            in1 => \N__33659\,
            in2 => \N__33441\,
            in3 => \N__33231\,
            lcout => \pwmWrite_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15684\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15675\,
            in2 => \N__32472\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_0\,
            carryout => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15666\,
            in2 => \N__32466\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_1\,
            carryout => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15651\,
            in2 => \N__32470\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_2\,
            carryout => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15783\,
            in2 => \N__32468\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_3\,
            carryout => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15771\,
            in2 => \N__32471\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_4\,
            carryout => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15759\,
            in2 => \N__32467\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_5\,
            carryout => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15747\,
            in2 => \N__32469\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_6\,
            carryout => \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.out_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__15725\,
            in1 => \N__16833\,
            in2 => \N__16999\,
            in3 => \N__15738\,
            lcout => \PWM1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38559\,
            ce => 'H',
            sr => \N__35719\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_13_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28723\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38552\,
            ce => \N__18233\,
            sr => \N__35727\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_5_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36367\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38552\,
            ce => \N__18233\,
            sr => \N__35727\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_8_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28992\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38552\,
            ce => \N__18233\,
            sr => \N__35727\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_9_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28576\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38552\,
            ce => \N__18233\,
            sr => \N__35727\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_12_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28870\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38552\,
            ce => \N__18233\,
            sr => \N__35727\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_6_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31114\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38552\,
            ce => \N__18233\,
            sr => \N__35727\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_4_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36513\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38552\,
            ce => \N__18233\,
            sr => \N__35727\
        );

    \PWMInstance0.periodCounter_RNIB5GO1_11_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15938\,
            in1 => \N__16904\,
            in2 => \N__17088\,
            in3 => \N__15983\,
            lcout => \PWMInstance0.un1_periodCounter12_1_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__16005\,
            in1 => \N__15807\,
            in2 => \N__15984\,
            in3 => \N__15813\,
            lcout => \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_2_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31603\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38548\,
            ce => \N__18235\,
            sr => \N__35738\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_3_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32082\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38548\,
            ce => \N__18235\,
            sr => \N__35738\
        );

    \PWMInstance0.periodCounter_RNIR3TO_14_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17147\,
            in2 => \_gnd_net_\,
            in3 => \N__16004\,
            lcout => OPEN,
            ltout => \PWMInstance0.un1_periodCounter12_1_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.periodCounter_RNIPQTQ1_10_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15960\,
            in1 => \N__17027\,
            in2 => \N__15798\,
            in3 => \N__17112\,
            lcout => \PWMInstance0.un1_periodCounter12_1_0_a2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__15795\,
            in1 => \N__15959\,
            in2 => \N__15939\,
            in3 => \N__15789\,
            lcout => \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.out_RNO_0_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15868\,
            in1 => \N__15900\,
            in2 => \N__15888\,
            in3 => \N__16062\,
            lcout => \PWMInstance0.un1_periodCounter12_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.clkCount_0_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__16874\,
            in1 => \N__15886\,
            in2 => \_gnd_net_\,
            in3 => \N__15869\,
            lcout => \PWMInstance0.clkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38545\,
            ce => 'H',
            sr => \N__35742\
        );

    \PWMInstance0.clkCount_1_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110001000"
        )
    port map (
            in0 => \N__16875\,
            in1 => \N__15887\,
            in2 => \_gnd_net_\,
            in3 => \N__15870\,
            lcout => \PWMInstance0.clkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38545\,
            ce => 'H',
            sr => \N__35742\
        );

    \PWMInstance0.periodCounter_RNI2BTO_16_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16061\,
            in2 => \_gnd_net_\,
            in3 => \N__17194\,
            lcout => \PWMInstance0.un1_periodCounter12_1_0_a2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.clkCount_RNIPL0S_0_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15899\,
            in1 => \N__15882\,
            in2 => \_gnd_net_\,
            in3 => \N__15867\,
            lcout => \PWMInstance0.periodCounter12\,
            ltout => \PWMInstance0.periodCounter12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.periodCounter_RNIM4RD2_15_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__17171\,
            in1 => \N__18007\,
            in2 => \N__15855\,
            in3 => \N__15852\,
            lcout => OPEN,
            ltout => \PWMInstance0.un1_periodCounter12_1_0_a2_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.periodCounter_RNI49PP7_10_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15846\,
            in1 => \N__18045\,
            in2 => \N__15840\,
            in3 => \N__15837\,
            lcout => \PWMInstance0.out_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.periodCounter_0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18034\,
            in2 => \N__15831\,
            in3 => \N__15830\,
            lcout => \PWMInstance0.periodCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_0\,
            clk => \N__38544\,
            ce => 'H',
            sr => \N__35303\
        );

    \PWMInstance0.periodCounter_1_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18011\,
            in2 => \_gnd_net_\,
            in3 => \N__15816\,
            lcout => \PWMInstance0.periodCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_0\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_1\,
            clk => \N__38544\,
            ce => 'H',
            sr => \N__35303\
        );

    \PWMInstance0.periodCounter_2_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16003\,
            in2 => \_gnd_net_\,
            in3 => \N__15987\,
            lcout => \PWMInstance0.periodCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_1\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_2\,
            clk => \N__38544\,
            ce => 'H',
            sr => \N__35303\
        );

    \PWMInstance0.periodCounter_3_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15979\,
            in2 => \_gnd_net_\,
            in3 => \N__15963\,
            lcout => \PWMInstance0.periodCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_2\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_3\,
            clk => \N__38544\,
            ce => 'H',
            sr => \N__35303\
        );

    \PWMInstance0.periodCounter_4_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15958\,
            in2 => \_gnd_net_\,
            in3 => \N__15942\,
            lcout => \PWMInstance0.periodCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_3\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_4\,
            clk => \N__38544\,
            ce => 'H',
            sr => \N__35303\
        );

    \PWMInstance0.periodCounter_5_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15934\,
            in2 => \_gnd_net_\,
            in3 => \N__15918\,
            lcout => \PWMInstance0.periodCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_4\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_5\,
            clk => \N__38544\,
            ce => 'H',
            sr => \N__35303\
        );

    \PWMInstance0.periodCounter_6_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18100\,
            in2 => \_gnd_net_\,
            in3 => \N__15915\,
            lcout => \PWMInstance0.periodCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_5\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_6\,
            clk => \N__38544\,
            ce => 'H',
            sr => \N__35303\
        );

    \PWMInstance0.periodCounter_7_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17284\,
            in1 => \N__17198\,
            in2 => \_gnd_net_\,
            in3 => \N__15912\,
            lcout => \PWMInstance0.periodCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_6\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_7\,
            clk => \N__38544\,
            ce => 'H',
            sr => \N__35303\
        );

    \PWMInstance0.periodCounter_8_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18133\,
            in2 => \_gnd_net_\,
            in3 => \N__15909\,
            lcout => \PWMInstance0.periodCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_8\,
            clk => \N__38543\,
            ce => 'H',
            sr => \N__35301\
        );

    \PWMInstance0.periodCounter_9_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16900\,
            in2 => \_gnd_net_\,
            in3 => \N__15906\,
            lcout => \PWMInstance0.periodCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_8\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_9\,
            clk => \N__38543\,
            ce => 'H',
            sr => \N__35301\
        );

    \PWMInstance0.periodCounter_10_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17110\,
            in2 => \_gnd_net_\,
            in3 => \N__15903\,
            lcout => \PWMInstance0.periodCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_9\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_10\,
            clk => \N__38543\,
            ce => 'H',
            sr => \N__35301\
        );

    \PWMInstance0.periodCounter_11_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17289\,
            in1 => \N__17080\,
            in2 => \_gnd_net_\,
            in3 => \N__16080\,
            lcout => \PWMInstance0.periodCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_10\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_11\,
            clk => \N__38543\,
            ce => 'H',
            sr => \N__35301\
        );

    \PWMInstance0.periodCounter_12_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17291\,
            in1 => \N__17026\,
            in2 => \_gnd_net_\,
            in3 => \N__16077\,
            lcout => \PWMInstance0.periodCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_11\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_12\,
            clk => \N__38543\,
            ce => 'H',
            sr => \N__35301\
        );

    \PWMInstance0.periodCounter_13_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17288\,
            in1 => \N__18067\,
            in2 => \_gnd_net_\,
            in3 => \N__16074\,
            lcout => \PWMInstance0.periodCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_12\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_13\,
            clk => \N__38543\,
            ce => 'H',
            sr => \N__35301\
        );

    \PWMInstance0.periodCounter_14_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17146\,
            in2 => \_gnd_net_\,
            in3 => \N__16071\,
            lcout => \PWMInstance0.periodCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_13\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_14\,
            clk => \N__38543\,
            ce => 'H',
            sr => \N__35301\
        );

    \PWMInstance0.periodCounter_15_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17170\,
            in2 => \_gnd_net_\,
            in3 => \N__16068\,
            lcout => \PWMInstance0.periodCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_periodCounter_2_cry_14\,
            carryout => \PWMInstance0.un1_periodCounter_2_cry_15\,
            clk => \N__38543\,
            ce => 'H',
            sr => \N__35301\
        );

    \PWMInstance0.periodCounter_16_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17290\,
            in1 => \N__16060\,
            in2 => \_gnd_net_\,
            in3 => \N__16065\,
            lcout => \PWMInstance0.periodCounterZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38541\,
            ce => 'H',
            sr => \N__35299\
        );

    \PWMInstance1.periodCounter_0_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16042\,
            in2 => \N__16596\,
            in3 => \N__16595\,
            lcout => \PWMInstance1.periodCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_0\,
            clk => \N__38678\,
            ce => 'H',
            sr => \N__35316\
        );

    \PWMInstance1.periodCounter_1_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16618\,
            in2 => \_gnd_net_\,
            in3 => \N__16026\,
            lcout => \PWMInstance1.periodCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_0\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_1\,
            clk => \N__38678\,
            ce => 'H',
            sr => \N__35316\
        );

    \PWMInstance1.periodCounter_2_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16023\,
            in2 => \_gnd_net_\,
            in3 => \N__16008\,
            lcout => \PWMInstance1.periodCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_1\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_2\,
            clk => \N__38678\,
            ce => 'H',
            sr => \N__35316\
        );

    \PWMInstance1.periodCounter_3_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16241\,
            in2 => \_gnd_net_\,
            in3 => \N__16224\,
            lcout => \PWMInstance1.periodCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_2\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_3\,
            clk => \N__38678\,
            ce => 'H',
            sr => \N__35316\
        );

    \PWMInstance1.periodCounter_4_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16221\,
            in2 => \_gnd_net_\,
            in3 => \N__16206\,
            lcout => \PWMInstance1.periodCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_3\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_4\,
            clk => \N__38678\,
            ce => 'H',
            sr => \N__35316\
        );

    \PWMInstance1.periodCounter_5_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16202\,
            in2 => \_gnd_net_\,
            in3 => \N__16185\,
            lcout => \PWMInstance1.periodCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_4\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_5\,
            clk => \N__38678\,
            ce => 'H',
            sr => \N__35316\
        );

    \PWMInstance1.periodCounter_6_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16172\,
            in2 => \_gnd_net_\,
            in3 => \N__16158\,
            lcout => \PWMInstance1.periodCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_5\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_6\,
            clk => \N__38678\,
            ce => 'H',
            sr => \N__35316\
        );

    \PWMInstance1.periodCounter_7_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17000\,
            in1 => \N__16678\,
            in2 => \_gnd_net_\,
            in3 => \N__16155\,
            lcout => \PWMInstance1.periodCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_6\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_7\,
            clk => \N__38678\,
            ce => 'H',
            sr => \N__35316\
        );

    \PWMInstance1.periodCounter_8_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16152\,
            in2 => \_gnd_net_\,
            in3 => \N__16134\,
            lcout => \PWMInstance1.periodCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_8\,
            clk => \N__38671\,
            ce => 'H',
            sr => \N__35315\
        );

    \PWMInstance1.periodCounter_9_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16130\,
            in2 => \_gnd_net_\,
            in3 => \N__16110\,
            lcout => \PWMInstance1.periodCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_8\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_9\,
            clk => \N__38671\,
            ce => 'H',
            sr => \N__35315\
        );

    \PWMInstance1.periodCounter_10_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16103\,
            in2 => \_gnd_net_\,
            in3 => \N__16083\,
            lcout => \PWMInstance1.periodCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_9\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_10\,
            clk => \N__38671\,
            ce => 'H',
            sr => \N__35315\
        );

    \PWMInstance1.periodCounter_11_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17002\,
            in1 => \N__16348\,
            in2 => \_gnd_net_\,
            in3 => \N__16326\,
            lcout => \PWMInstance1.periodCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_10\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_11\,
            clk => \N__38671\,
            ce => 'H',
            sr => \N__35315\
        );

    \PWMInstance1.periodCounter_12_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17004\,
            in1 => \N__16322\,
            in2 => \_gnd_net_\,
            in3 => \N__16302\,
            lcout => \PWMInstance1.periodCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_11\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_12\,
            clk => \N__38671\,
            ce => 'H',
            sr => \N__35315\
        );

    \PWMInstance1.periodCounter_13_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17003\,
            in1 => \N__16294\,
            in2 => \_gnd_net_\,
            in3 => \N__16275\,
            lcout => \PWMInstance1.periodCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_12\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_13\,
            clk => \N__38671\,
            ce => 'H',
            sr => \N__35315\
        );

    \PWMInstance1.periodCounter_14_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16271\,
            in2 => \_gnd_net_\,
            in3 => \N__16251\,
            lcout => \PWMInstance1.periodCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_13\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_14\,
            clk => \N__38671\,
            ce => 'H',
            sr => \N__35315\
        );

    \PWMInstance1.periodCounter_15_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16648\,
            in2 => \_gnd_net_\,
            in3 => \N__16248\,
            lcout => \PWMInstance1.periodCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \PWMInstance1.un1_periodCounter_2_cry_14\,
            carryout => \PWMInstance1.un1_periodCounter_2_cry_15\,
            clk => \N__38671\,
            ce => 'H',
            sr => \N__35315\
        );

    \PWMInstance1.periodCounter_16_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17001\,
            in1 => \N__16702\,
            in2 => \_gnd_net_\,
            in3 => \N__16245\,
            lcout => \PWMInstance1.periodCounterZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38659\,
            ce => 'H',
            sr => \N__35313\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17907\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16962\,
            in2 => \N__32592\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_0\,
            carryout => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19272\,
            in2 => \N__32586\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_1\,
            carryout => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17883\,
            in2 => \N__32590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_2\,
            carryout => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16416\,
            in2 => \N__32588\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_3\,
            carryout => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19143\,
            in2 => \N__32591\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_4\,
            carryout => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17220\,
            in2 => \N__32587\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_5\,
            carryout => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16932\,
            in2 => \N__32589\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_6\,
            carryout => \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.out_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__16385\,
            in1 => \N__19122\,
            in2 => \N__19461\,
            in3 => \N__16404\,
            lcout => \PWM5_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38639\,
            ce => 'H',
            sr => \N__35682\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_12_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28875\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38628\,
            ce => \N__16803\,
            sr => \N__35685\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_10_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36168\,
            lcout => \PWMInstance1.PWMPulseWidthCountZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38628\,
            ce => \N__16803\,
            sr => \N__35685\
        );

    \QuadInstance2.Quad_9_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28577\,
            in2 => \N__16359\,
            in3 => \N__22142\,
            lcout => \dataRead2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38617\,
            ce => 'H',
            sr => \N__35691\
        );

    \QuadInstance2.Quad_10_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22139\,
            in1 => \N__36160\,
            in2 => \_gnd_net_\,
            in3 => \N__16434\,
            lcout => \dataRead2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38617\,
            ce => 'H',
            sr => \N__35691\
        );

    \QuadInstance7.Quad_11_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__36011\,
            in1 => \_gnd_net_\,
            in2 => \N__26037\,
            in3 => \N__17727\,
            lcout => \dataRead7_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38617\,
            ce => 'H',
            sr => \N__35691\
        );

    \QuadInstance4.Quad_9_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28578\,
            in1 => \N__29662\,
            in2 => \_gnd_net_\,
            in3 => \N__25050\,
            lcout => \dataRead4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38617\,
            ce => 'H',
            sr => \N__35691\
        );

    \QuadInstance2.Quad_14_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34403\,
            in1 => \N__22141\,
            in2 => \_gnd_net_\,
            in3 => \N__16428\,
            lcout => \dataRead2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38617\,
            ce => 'H',
            sr => \N__35691\
        );

    \QuadInstance1.Quad_2_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31593\,
            in1 => \N__24086\,
            in2 => \_gnd_net_\,
            in3 => \N__21633\,
            lcout => \dataRead1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38617\,
            ce => 'H',
            sr => \N__35691\
        );

    \QuadInstance7.Quad_12_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26004\,
            in1 => \N__28866\,
            in2 => \_gnd_net_\,
            in3 => \N__17706\,
            lcout => \dataRead7_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38617\,
            ce => 'H',
            sr => \N__35691\
        );

    \QuadInstance2.Quad_12_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22140\,
            in1 => \_gnd_net_\,
            in2 => \N__28874\,
            in3 => \N__16422\,
            lcout => \dataRead2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38617\,
            ce => 'H',
            sr => \N__35691\
        );

    \quadWrite_2_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33225\,
            in1 => \N__33848\,
            in2 => \N__33450\,
            in3 => \N__33652\,
            lcout => \quadWriteZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIB8VV2_4_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__21465\,
            in1 => \N__25920\,
            in2 => \N__21800\,
            in3 => \N__16512\,
            lcout => \QuadInstance7.Quad_RNIB8VV2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quadWrite_7_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33847\,
            in1 => \N__33651\,
            in2 => \N__33451\,
            in3 => \N__23458\,
            lcout => \quadWriteZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIA7VV2_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__27842\,
            in1 => \N__25919\,
            in2 => \N__21799\,
            in3 => \N__16510\,
            lcout => \QuadInstance7.Quad_RNIA7VV2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIDAVV2_6_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__16513\,
            in1 => \N__27704\,
            in2 => \N__25971\,
            in3 => \N__21781\,
            lcout => \QuadInstance7.Quad_RNIDAVV2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIEBVV2_7_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__26271\,
            in1 => \N__25927\,
            in2 => \N__21801\,
            in3 => \N__16514\,
            lcout => \QuadInstance7.Quad_RNIEBVV2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIC9VV2_5_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__16511\,
            in1 => \N__36746\,
            in2 => \N__25970\,
            in3 => \N__21777\,
            lcout => \QuadInstance7.Quad_RNIC9VV2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIOIKU2_10_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001100"
        )
    port map (
            in0 => \N__34650\,
            in1 => \N__21787\,
            in2 => \N__25973\,
            in3 => \N__16508\,
            lcout => \QuadInstance7.Quad_RNIOIKU2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.delayedCh_B_RNI2N241_2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34470\,
            in1 => \N__16841\,
            in2 => \_gnd_net_\,
            in3 => \N__16462\,
            lcout => \QuadInstance7.un1_count_enable_i_a2_0_1\,
            ltout => \QuadInstance7.un1_count_enable_i_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNI96VV2_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__30386\,
            in1 => \N__25918\,
            in2 => \N__16440\,
            in3 => \N__21782\,
            lcout => \QuadInstance7.Quad_RNI96VV2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.delayedCh_A_RNI8MRP1_2_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16853\,
            in1 => \N__16463\,
            in2 => \N__16449\,
            in3 => \N__16842\,
            lcout => \QuadInstance7.count_enable\,
            ltout => \QuadInstance7.count_enable_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNI85VV2_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__25841\,
            in1 => \N__25917\,
            in2 => \N__16437\,
            in3 => \N__16505\,
            lcout => \QuadInstance7.Quad_RNI85VV2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIFCVV2_8_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011010000"
        )
    port map (
            in0 => \N__16506\,
            in1 => \N__25928\,
            in2 => \N__21802\,
            in3 => \N__37613\,
            lcout => \QuadInstance7.Quad_RNIFCVV2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIGDVV2_9_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001100"
        )
    port map (
            in0 => \N__25392\,
            in1 => \N__21786\,
            in2 => \N__25972\,
            in3 => \N__16507\,
            lcout => \QuadInstance7.Quad_RNIGDVV2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIRLKU2_13_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011010000"
        )
    port map (
            in0 => \N__16509\,
            in1 => \N__25935\,
            in2 => \N__21803\,
            in3 => \N__26112\,
            lcout => \QuadInstance7.Quad_RNIRLKU2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNISMKU2_14_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__16521\,
            in1 => \N__25976\,
            in2 => \N__20283\,
            in3 => \N__21794\,
            lcout => \QuadInstance7.Quad_RNISMKU2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.delayedCh_B_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17418\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance7.delayedCh_BZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIPJKU2_11_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__20877\,
            in1 => \N__25974\,
            in2 => \N__16523\,
            in3 => \N__21792\,
            lcout => \QuadInstance7.Quad_RNIPJKU2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.delayedCh_A_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29694\,
            lcout => \QuadInstance7.delayedCh_AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNIQKKU2_12_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__22262\,
            in1 => \N__25975\,
            in2 => \N__16524\,
            in3 => \N__21793\,
            lcout => \QuadInstance7.Quad_RNIQKKU2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__23451\,
            in1 => \N__33830\,
            in2 => \N__33442\,
            in3 => \N__33666\,
            lcout => \pwmWriteZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.delayedCh_A_2_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16464\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance7.delayedCh_AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.delayedCh_B_2_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16854\,
            lcout => \QuadInstance7.delayedCh_BZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.out_RNO_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__17823\,
            in1 => \N__16735\,
            in2 => \N__16707\,
            in3 => \N__16720\,
            lcout => \PWMInstance1.un1_periodCounter12_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.clkCount_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000101"
        )
    port map (
            in0 => \N__16721\,
            in1 => \_gnd_net_\,
            in2 => \N__16742\,
            in3 => \N__16754\,
            lcout => \PWMInstance1.clkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38576\,
            ce => 'H',
            sr => \N__35720\
        );

    \PWMInstance1.PWMPulseWidthCount_esr_ctle_15_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__16753\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35825\,
            lcout => \PWMInstance1.pwmWrite_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.clkCount_1_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000001010"
        )
    port map (
            in0 => \N__16722\,
            in1 => \_gnd_net_\,
            in2 => \N__16743\,
            in3 => \N__16755\,
            lcout => \PWMInstance1.clkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38576\,
            ce => 'H',
            sr => \N__35720\
        );

    \PWMInstance1.clkCount_RNISE5O_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__17822\,
            in1 => \N__16734\,
            in2 => \_gnd_net_\,
            in3 => \N__16719\,
            lcout => \PWMInstance1.periodCounter12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.periodCounter_RNI4EVP_16_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16703\,
            in2 => \_gnd_net_\,
            in3 => \N__16686\,
            lcout => OPEN,
            ltout => \PWMInstance1.un1_periodCounter12_1_0_a2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.periodCounter_RNIT34C2_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__16655\,
            in1 => \N__16626\,
            in2 => \N__16599\,
            in3 => \N__16580\,
            lcout => OPEN,
            ltout => \PWMInstance1.un1_periodCounter12_1_0_a2_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance1.periodCounter_RNIOA6I7_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16569\,
            in1 => \N__16554\,
            in2 => \N__16542\,
            in3 => \N__16539\,
            lcout => \PWMInstance1.out_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__16947\,
            in1 => \N__16953\,
            in2 => \N__19346\,
            in3 => \N__19256\,
            lcout => \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_2_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31591\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38566\,
            ce => \N__19635\,
            sr => \N__35728\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32085\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38566\,
            ce => \N__19635\,
            sr => \N__35728\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__16941\,
            in1 => \N__16920\,
            in2 => \N__19524\,
            in3 => \N__19238\,
            lcout => \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_15_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31871\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38566\,
            ce => \N__19635\,
            sr => \N__35728\
        );

    \pwmWrite_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__33849\,
            in1 => \N__33672\,
            in2 => \N__33452\,
            in3 => \N__33224\,
            lcout => \pwmWriteZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__18140\,
            in1 => \N__16914\,
            in2 => \N__16908\,
            in3 => \N__16881\,
            lcout => \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_ctle_15_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__35826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16865\,
            lcout => \PWMInstance0.pwmWrite_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__18210\,
            in1 => \N__17232\,
            in2 => \N__18177\,
            in3 => \N__19220\,
            lcout => \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__18261\,
            in1 => \N__17208\,
            in2 => \N__18111\,
            in3 => \N__17202\,
            lcout => \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__17118\,
            in1 => \N__17124\,
            in2 => \N__17178\,
            in3 => \N__17151\,
            lcout => \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_14_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34378\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38553\,
            ce => \N__18234\,
            sr => \N__35743\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_15_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31878\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38553\,
            ce => \N__18234\,
            sr => \N__35743\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__17111\,
            in1 => \N__17046\,
            in2 => \N__17087\,
            in3 => \N__17058\,
            lcout => \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_11_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35998\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38553\,
            ce => \N__18234\,
            sr => \N__35743\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__17040\,
            in1 => \N__17034\,
            in2 => \N__18077\,
            in3 => \N__17028\,
            lcout => \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17988\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17346\,
            in2 => \N__32572\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_0\,
            carryout => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17340\,
            in2 => \N__32566\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_1\,
            carryout => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17334\,
            in2 => \N__32570\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_2\,
            carryout => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17325\,
            in2 => \N__32568\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_3\,
            carryout => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17316\,
            in2 => \N__32571\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_4\,
            carryout => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17310\,
            in2 => \N__32567\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_5\,
            carryout => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17304\,
            in2 => \N__32569\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_6\,
            carryout => \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.out_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__17243\,
            in1 => \N__17298\,
            in2 => \N__17292\,
            in3 => \N__17253\,
            lcout => \PWM0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38546\,
            ce => 'H',
            sr => \N__35755\
        );

    \QuadInstance7.delayedCh_B_0_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17436\,
            lcout => \QuadInstance7.delayedCh_BZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38542\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM0_obufLegalizeSB_DFF_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM0_obufLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM1_obufLegalizeSB_DFF_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM1_obufLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM6_obufLegalizeSB_DFF_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM6_obufLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM7_obufLegalizeSB_DFF_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM7_obufLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.delayedCh_B_0_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17385\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance3.delayedCh_BZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_4_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36521\,
            in1 => \N__22171\,
            in2 => \_gnd_net_\,
            in3 => \N__17376\,
            lcout => \dataRead2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38672\,
            ce => 'H',
            sr => \N__35681\
        );

    \QuadInstance5.delayedCh_A_1_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17352\,
            lcout => \QuadInstance5.delayedCh_AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.delayedCh_A_0_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17364\,
            lcout => \QuadInstance5.delayedCh_AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNI07LI2_9_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__25514\,
            in1 => \N__25727\,
            in2 => \N__17500\,
            in3 => \N__18368\,
            lcout => \QuadInstance5.Quad_RNI07LI2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.delayedCh_B_RNIUQSQ_2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34500\,
            in1 => \N__18407\,
            in2 => \_gnd_net_\,
            in3 => \N__18433\,
            lcout => \QuadInstance5.un1_count_enable_i_a2_0_1\,
            ltout => \QuadInstance5.un1_count_enable_i_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIPVKI2_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__30530\,
            in1 => \N__25723\,
            in2 => \N__17439\,
            in3 => \N__18360\,
            lcout => \QuadInstance5.Quad_RNIPVKI2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIQ0LI2_3_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__27918\,
            in1 => \N__25724\,
            in2 => \N__17499\,
            in3 => \N__18364\,
            lcout => \QuadInstance5.Quad_RNIQ0LI2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIR1LI2_4_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__25725\,
            in1 => \N__21326\,
            in2 => \N__18382\,
            in3 => \N__17478\,
            lcout => \QuadInstance5.Quad_RNIR1LI2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIS2LI2_5_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__25726\,
            in1 => \N__36871\,
            in2 => \N__18383\,
            in3 => \N__17482\,
            lcout => \QuadInstance5.Quad_RNIS2LI2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNI8AQ82_10_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__25722\,
            in1 => \N__17486\,
            in2 => \N__35024\,
            in3 => \N__18358\,
            lcout => \QuadInstance5.Quad_RNI8AQ82Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNI9BQ82_11_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001010"
        )
    port map (
            in0 => \N__18359\,
            in1 => \N__25721\,
            in2 => \N__17501\,
            in3 => \N__20112\,
            lcout => \QuadInstance5.Quad_RNI9BQ82Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quadWrite_5_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33827\,
            in1 => \N__33639\,
            in2 => \N__33466\,
            in3 => \N__23459\,
            lcout => \quadWriteZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIT3LI2_6_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__25281\,
            in1 => \N__25716\,
            in2 => \N__18380\,
            in3 => \N__17476\,
            lcout => \QuadInstance5.Quad_RNIT3LI2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIU4LI2_7_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__17475\,
            in1 => \N__25607\,
            in2 => \N__25757\,
            in3 => \N__18351\,
            lcout => \QuadInstance5.Quad_RNIU4LI2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIV5LI2_8_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__36984\,
            in1 => \N__25720\,
            in2 => \N__18381\,
            in3 => \N__17477\,
            lcout => \QuadInstance5.Quad_RNIV5LI2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_RNIJ03G2_13_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__19974\,
            in1 => \N__22143\,
            in2 => \N__17601\,
            in3 => \N__18530\,
            lcout => \QuadInstance2.Quad_RNIJ03G2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIOUKI2_1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__23858\,
            in1 => \N__25715\,
            in2 => \N__18379\,
            in3 => \N__17474\,
            lcout => \QuadInstance5.Quad_RNIOUKI2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIACQ82_12_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__25728\,
            in1 => \N__17503\,
            in2 => \N__22385\,
            in3 => \N__18387\,
            lcout => \QuadInstance5.Quad_RNIACQ82Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNIBDQ82_13_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010000"
        )
    port map (
            in0 => \N__17502\,
            in1 => \N__20008\,
            in2 => \N__18392\,
            in3 => \N__25729\,
            lcout => \QuadInstance5.Quad_RNIBDQ82Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNICEQ82_14_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__25730\,
            in1 => \N__18388\,
            in2 => \N__28222\,
            in3 => \N__17504\,
            lcout => \QuadInstance5.Quad_RNICEQ82Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_15_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010011100"
        )
    port map (
            in0 => \N__17505\,
            in1 => \N__24242\,
            in2 => \N__18393\,
            in3 => \N__25731\,
            lcout => \QuadInstance5.un1_Quad_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_12_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25732\,
            in1 => \N__28847\,
            in2 => \_gnd_net_\,
            in3 => \N__18543\,
            lcout => \dataRead5_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38629\,
            ce => 'H',
            sr => \N__35698\
        );

    \QuadInstance5.Quad_13_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28719\,
            in1 => \N__25734\,
            in2 => \_gnd_net_\,
            in3 => \N__18705\,
            lcout => \dataRead5_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38629\,
            ce => 'H',
            sr => \N__35698\
        );

    \QuadInstance5.Quad_14_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25733\,
            in1 => \N__34402\,
            in2 => \_gnd_net_\,
            in3 => \N__18690\,
            lcout => \dataRead5_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38629\,
            ce => 'H',
            sr => \N__35698\
        );

    \QuadInstance5.Quad_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31248\,
            in1 => \N__18300\,
            in2 => \_gnd_net_\,
            in3 => \N__25735\,
            lcout => \dataRead5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38629\,
            ce => 'H',
            sr => \N__35698\
        );

    \QuadInstance7.un1_Quad_cry_0_c_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21791\,
            in2 => \N__30776\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \QuadInstance7.un1_Quad_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25842\,
            in2 => \N__17673\,
            in3 => \N__17664\,
            lcout => \QuadInstance7.Quad_RNO_0_6_1\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_0\,
            carryout => \QuadInstance7.un1_Quad_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30379\,
            in2 => \N__17661\,
            in3 => \N__17652\,
            lcout => \QuadInstance7.Quad_RNO_0_7_2\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_1\,
            carryout => \QuadInstance7.un1_Quad_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27841\,
            in2 => \N__17649\,
            in3 => \N__17640\,
            lcout => \QuadInstance7.Quad_RNO_0_7_3\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_2\,
            carryout => \QuadInstance7.un1_Quad_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_4_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21464\,
            in2 => \N__17637\,
            in3 => \N__17628\,
            lcout => \QuadInstance7.Quad_RNO_0_7_4\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_3\,
            carryout => \QuadInstance7.un1_Quad_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_5_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36739\,
            in2 => \N__17625\,
            in3 => \N__17616\,
            lcout => \QuadInstance7.Quad_RNO_0_7_5\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_4\,
            carryout => \QuadInstance7.un1_Quad_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_6_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27700\,
            in2 => \N__17613\,
            in3 => \N__17604\,
            lcout => \QuadInstance7.Quad_RNO_0_7_6\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_5\,
            carryout => \QuadInstance7.un1_Quad_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_7_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26257\,
            in2 => \N__17784\,
            in3 => \N__17775\,
            lcout => \QuadInstance7.Quad_RNO_0_7_7\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_6\,
            carryout => \QuadInstance7.un1_Quad_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_8_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37612\,
            in2 => \N__17772\,
            in3 => \N__17763\,
            lcout => \QuadInstance7.Quad_RNO_0_7_8\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \QuadInstance7.un1_Quad_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_9_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25387\,
            in2 => \N__17760\,
            in3 => \N__17751\,
            lcout => \QuadInstance7.Quad_RNO_0_7_9\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_8\,
            carryout => \QuadInstance7.un1_Quad_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_10_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34645\,
            in2 => \N__17748\,
            in3 => \N__17739\,
            lcout => \QuadInstance7.Quad_RNO_0_7_10\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_9\,
            carryout => \QuadInstance7.un1_Quad_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_11_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20875\,
            in2 => \N__17736\,
            in3 => \N__17718\,
            lcout => \QuadInstance7.Quad_RNO_0_7_11\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_10\,
            carryout => \QuadInstance7.un1_Quad_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_12_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22252\,
            in2 => \N__17715\,
            in3 => \N__17697\,
            lcout => \QuadInstance7.Quad_RNO_0_7_12\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_11\,
            carryout => \QuadInstance7.un1_Quad_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_13_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26108\,
            in2 => \N__17694\,
            in3 => \N__17685\,
            lcout => \QuadInstance7.Quad_RNO_0_7_13\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_12\,
            carryout => \QuadInstance7.un1_Quad_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_RNO_0_14_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17682\,
            in2 => \N__20282\,
            in3 => \N__17676\,
            lcout => \QuadInstance7.Quad_RNO_0_7_14\,
            ltout => OPEN,
            carryin => \QuadInstance7.un1_Quad_cry_13\,
            carryout => \QuadInstance7.un1_Quad_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance7.Quad_15_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__17835\,
            in1 => \N__25969\,
            in2 => \N__31909\,
            in3 => \N__17826\,
            lcout => \dataRead7_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38608\,
            ce => 'H',
            sr => \N__35709\
        );

    \QuadInstance3.Quad_RNIQ30J1_12_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__21928\,
            in1 => \N__19035\,
            in2 => \N__22332\,
            in3 => \N__18947\,
            lcout => \QuadInstance3.Quad_RNIQ30J1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIAQAL1_3_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__24375\,
            in1 => \N__21922\,
            in2 => \N__18971\,
            in3 => \N__19024\,
            lcout => \QuadInstance3.Quad_RNIAQAL1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIDTAL1_6_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__19025\,
            in1 => \N__28265\,
            in2 => \N__21969\,
            in3 => \N__18945\,
            lcout => \QuadInstance3.Quad_RNIDTAL1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNICSAL1_5_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__23745\,
            in1 => \N__21923\,
            in2 => \N__18972\,
            in3 => \N__19026\,
            lcout => \QuadInstance3.Quad_RNICSAL1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIR40J1_13_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__21929\,
            in1 => \N__19039\,
            in2 => \N__19938\,
            in3 => \N__18948\,
            lcout => \QuadInstance3.Quad_RNIR40J1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIP20J1_11_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001010"
        )
    port map (
            in0 => \N__18946\,
            in1 => \N__21927\,
            in2 => \N__19041\,
            in3 => \N__22422\,
            lcout => \QuadInstance3.Quad_RNIP20J1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_fast_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__23450\,
            in1 => \N__33367\,
            in2 => \N__33671\,
            in3 => \N__33829\,
            lcout => \pwmWrite_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_7_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__33828\,
            in1 => \N__33662\,
            in2 => \N__33432\,
            in3 => \N__23449\,
            lcout => \pwmWriteZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.periodCounter_RNIUTF81_13_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__17855\,
            in1 => \N__18173\,
            in2 => \N__17967\,
            in3 => \N__17943\,
            lcout => \PWMInstance5.un1_periodCounter12_1_0_a2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__17889\,
            in1 => \N__17854\,
            in2 => \N__19503\,
            in3 => \N__17895\,
            lcout => \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31374\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38588\,
            ce => \N__19639\,
            sr => \N__35729\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31239\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38588\,
            ce => \N__19639\,
            sr => \N__35729\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__17962\,
            in1 => \N__17871\,
            in2 => \N__17865\,
            in3 => \N__19297\,
            lcout => \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_6_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31087\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38588\,
            ce => \N__19639\,
            sr => \N__35729\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_7_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29425\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38588\,
            ce => \N__19639\,
            sr => \N__35729\
        );

    \PWMInstance5.periodCounter_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17856\,
            in2 => \N__19539\,
            in3 => \N__19538\,
            lcout => \PWMInstance5.periodCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_0\,
            clk => \N__38577\,
            ce => 'H',
            sr => \N__35307\
        );

    \PWMInstance5.periodCounter_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19502\,
            in2 => \_gnd_net_\,
            in3 => \N__17841\,
            lcout => \PWMInstance5.periodCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_0\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_1\,
            clk => \N__38577\,
            ce => 'H',
            sr => \N__35307\
        );

    \PWMInstance5.periodCounter_2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19257\,
            in2 => \_gnd_net_\,
            in3 => \N__17838\,
            lcout => \PWMInstance5.periodCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_1\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_2\,
            clk => \N__38577\,
            ce => 'H',
            sr => \N__35307\
        );

    \PWMInstance5.periodCounter_3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19345\,
            in2 => \_gnd_net_\,
            in3 => \N__17976\,
            lcout => \PWMInstance5.periodCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_2\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_3\,
            clk => \N__38577\,
            ce => 'H',
            sr => \N__35307\
        );

    \PWMInstance5.periodCounter_4_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19200\,
            in2 => \_gnd_net_\,
            in3 => \N__17973\,
            lcout => \PWMInstance5.periodCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_3\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_4\,
            clk => \N__38577\,
            ce => 'H',
            sr => \N__35307\
        );

    \PWMInstance5.periodCounter_5_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19393\,
            in2 => \_gnd_net_\,
            in3 => \N__17970\,
            lcout => \PWMInstance5.periodCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_4\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_5\,
            clk => \N__38577\,
            ce => 'H',
            sr => \N__35307\
        );

    \PWMInstance5.periodCounter_6_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17966\,
            in2 => \_gnd_net_\,
            in3 => \N__17949\,
            lcout => \PWMInstance5.periodCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_5\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_6\,
            clk => \N__38577\,
            ce => 'H',
            sr => \N__35307\
        );

    \PWMInstance5.periodCounter_7_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19451\,
            in1 => \N__19298\,
            in2 => \_gnd_net_\,
            in3 => \N__17946\,
            lcout => \PWMInstance5.periodCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_6\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_7\,
            clk => \N__38577\,
            ce => 'H',
            sr => \N__35307\
        );

    \PWMInstance5.periodCounter_8_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17941\,
            in2 => \_gnd_net_\,
            in3 => \N__17919\,
            lcout => \PWMInstance5.periodCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_8\,
            clk => \N__38567\,
            ce => 'H',
            sr => \N__35306\
        );

    \PWMInstance5.periodCounter_9_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19415\,
            in2 => \_gnd_net_\,
            in3 => \N__17916\,
            lcout => \PWMInstance5.periodCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_8\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_9\,
            clk => \N__38567\,
            ce => 'H',
            sr => \N__35306\
        );

    \PWMInstance5.periodCounter_10_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19173\,
            in2 => \_gnd_net_\,
            in3 => \N__17913\,
            lcout => \PWMInstance5.periodCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_9\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_10\,
            clk => \N__38567\,
            ce => 'H',
            sr => \N__35306\
        );

    \PWMInstance5.periodCounter_11_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19453\,
            in1 => \N__19369\,
            in2 => \_gnd_net_\,
            in3 => \N__17910\,
            lcout => \PWMInstance5.periodCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_10\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_11\,
            clk => \N__38567\,
            ce => 'H',
            sr => \N__35306\
        );

    \PWMInstance5.periodCounter_12_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19450\,
            in1 => \N__19221\,
            in2 => \_gnd_net_\,
            in3 => \N__18180\,
            lcout => \PWMInstance5.periodCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_11\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_12\,
            clk => \N__38567\,
            ce => 'H',
            sr => \N__35306\
        );

    \PWMInstance5.periodCounter_13_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19454\,
            in1 => \N__18172\,
            in2 => \_gnd_net_\,
            in3 => \N__18153\,
            lcout => \PWMInstance5.periodCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_12\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_13\,
            clk => \N__38567\,
            ce => 'H',
            sr => \N__35306\
        );

    \PWMInstance5.periodCounter_14_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19239\,
            in2 => \_gnd_net_\,
            in3 => \N__18150\,
            lcout => \PWMInstance5.periodCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_13\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_14\,
            clk => \N__38567\,
            ce => 'H',
            sr => \N__35306\
        );

    \PWMInstance5.periodCounter_15_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19523\,
            in2 => \_gnd_net_\,
            in3 => \N__18147\,
            lcout => \PWMInstance5.periodCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \PWMInstance5.un1_periodCounter_2_cry_14\,
            carryout => \PWMInstance5.un1_periodCounter_2_cry_15\,
            clk => \N__38567\,
            ce => 'H',
            sr => \N__35306\
        );

    \PWMInstance5.periodCounter_16_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19452\,
            in1 => \N__19317\,
            in2 => \_gnd_net_\,
            in3 => \N__18144\,
            lcout => \PWMInstance5.periodCounterZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38561\,
            ce => 'H',
            sr => \N__35304\
        );

    \PWMInstance0.periodCounter_RNIA4GO1_13_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__18141\,
            in1 => \N__18110\,
            in2 => \N__18078\,
            in3 => \N__18036\,
            lcout => \PWMInstance0.un1_periodCounter12_1_0_a2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__18035\,
            in1 => \N__18267\,
            in2 => \N__18015\,
            in3 => \N__17982\,
            lcout => \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31422\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38554\,
            ce => \N__18248\,
            sr => \N__35756\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_1_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31264\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38554\,
            ce => \N__18248\,
            sr => \N__35756\
        );

    \PWMInstance0.PWMPulseWidthCount_esr_7_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29456\,
            lcout => \PWMInstance0.PWMPulseWidthCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38554\,
            ce => \N__18248\,
            sr => \N__35756\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_13_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28726\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38549\,
            ce => \N__19649\,
            sr => \N__35759\
        );

    \QuadInstance5.delayedCh_B_0_LC_10_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18201\,
            lcout => \QuadInstance5.delayedCh_BZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.delayedCh_A_2_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18435\,
            lcout => \QuadInstance5.delayedCh_AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.delayedCh_B_1_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18189\,
            lcout => \QuadInstance5.delayedCh_BZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.delayedCh_B_2_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18447\,
            lcout => \QuadInstance5.delayedCh_BZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_15_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111110000"
        )
    port map (
            in0 => \N__29663\,
            in1 => \N__27354\,
            in2 => \N__25224\,
            in3 => \N__27452\,
            lcout => \QuadInstance4.un1_Quad_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_0_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001100110"
        )
    port map (
            in0 => \N__27453\,
            in1 => \N__30268\,
            in2 => \N__31440\,
            in3 => \N__29664\,
            lcout => \dataRead4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38649\,
            ce => 'H',
            sr => \N__35689\
        );

    \QuadInstance0.Quad_0_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__30299\,
            in1 => \N__33127\,
            in2 => \N__31438\,
            in3 => \N__34089\,
            lcout => \dataRead0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38649\,
            ce => 'H',
            sr => \N__35689\
        );

    \QuadInstance2.Quad_0_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011000000110"
        )
    port map (
            in0 => \N__18534\,
            in1 => \N__30838\,
            in2 => \N__22190\,
            in3 => \N__31429\,
            lcout => \dataRead2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38649\,
            ce => 'H',
            sr => \N__35689\
        );

    \QuadInstance5.delayedCh_A_RNI0UF71_2_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18446\,
            in1 => \N__18434\,
            in2 => \N__18417\,
            in3 => \N__18408\,
            lcout => \QuadInstance5.count_enable\,
            ltout => \QuadInstance5.count_enable_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_0_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__25778\,
            in1 => \N__30907\,
            in2 => \N__18396\,
            in3 => \N__31430\,
            lcout => \dataRead5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38649\,
            ce => 'H',
            sr => \N__35689\
        );

    \QuadInstance3.Quad_0_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__22008\,
            in1 => \N__30877\,
            in2 => \N__31439\,
            in3 => \N__18978\,
            lcout => \dataRead3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38649\,
            ce => 'H',
            sr => \N__35689\
        );

    \QuadInstance5.un1_Quad_cry_0_c_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18369\,
            in2 => \N__30908\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_6_0_\,
            carryout => \QuadInstance5.un1_Quad_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_1_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23854\,
            in2 => \N__18309\,
            in3 => \N__18294\,
            lcout => \QuadInstance5.Quad_RNO_0_4_1\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_0\,
            carryout => \QuadInstance5.un1_Quad_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30526\,
            in2 => \N__18291\,
            in3 => \N__18282\,
            lcout => \QuadInstance5.Quad_RNO_0_5_2\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_1\,
            carryout => \QuadInstance5.un1_Quad_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_3_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27917\,
            in2 => \N__18279\,
            in3 => \N__18270\,
            lcout => \QuadInstance5.Quad_RNO_0_5_3\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_2\,
            carryout => \QuadInstance5.un1_Quad_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_4_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21316\,
            in2 => \N__18648\,
            in3 => \N__18639\,
            lcout => \QuadInstance5.Quad_RNO_0_5_4\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_3\,
            carryout => \QuadInstance5.un1_Quad_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_5_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36872\,
            in2 => \N__18636\,
            in3 => \N__18627\,
            lcout => \QuadInstance5.Quad_RNO_0_5_5\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_4\,
            carryout => \QuadInstance5.un1_Quad_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_6_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25267\,
            in2 => \N__18624\,
            in3 => \N__18615\,
            lcout => \QuadInstance5.Quad_RNO_0_5_6\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_5\,
            carryout => \QuadInstance5.un1_Quad_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_7_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18612\,
            in2 => \N__25597\,
            in3 => \N__18606\,
            lcout => \QuadInstance5.Quad_RNO_0_5_7\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_6\,
            carryout => \QuadInstance5.un1_Quad_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_8_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36973\,
            in2 => \N__18603\,
            in3 => \N__18594\,
            lcout => \QuadInstance5.Quad_RNO_0_5_8\,
            ltout => OPEN,
            carryin => \bfn_10_7_0_\,
            carryout => \QuadInstance5.un1_Quad_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_9_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25507\,
            in2 => \N__18591\,
            in3 => \N__18579\,
            lcout => \QuadInstance5.Quad_RNO_0_5_9\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_8\,
            carryout => \QuadInstance5.un1_Quad_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_10_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35008\,
            in2 => \N__18576\,
            in3 => \N__18567\,
            lcout => \QuadInstance5.Quad_RNO_0_5_10\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_9\,
            carryout => \QuadInstance5.un1_Quad_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_11_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20101\,
            in2 => \N__18564\,
            in3 => \N__18555\,
            lcout => \QuadInstance5.Quad_RNO_0_5_11\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_10\,
            carryout => \QuadInstance5.un1_Quad_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_12_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22378\,
            in2 => \N__18552\,
            in3 => \N__18537\,
            lcout => \QuadInstance5.Quad_RNO_0_5_12\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_11\,
            carryout => \QuadInstance5.un1_Quad_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_13_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18711\,
            in2 => \N__20012\,
            in3 => \N__18699\,
            lcout => \QuadInstance5.Quad_RNO_0_5_13\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_12\,
            carryout => \QuadInstance5.un1_Quad_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_RNO_0_14_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18696\,
            in2 => \N__28226\,
            in3 => \N__18684\,
            lcout => \QuadInstance5.Quad_RNO_0_5_14\,
            ltout => OPEN,
            carryin => \QuadInstance5.un1_Quad_cry_13\,
            carryout => \QuadInstance5.un1_Quad_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance5.Quad_15_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__18681\,
            in1 => \N__25756\,
            in2 => \N__31919\,
            in3 => \N__18675\,
            lcout => \dataRead5_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38630\,
            ce => 'H',
            sr => \N__35699\
        );

    \QuadInstance3.un1_Quad_cry_0_c_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18976\,
            in2 => \N__30878\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_8_0_\,
            carryout => \QuadInstance3.un1_Quad_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23807\,
            in2 => \N__18843\,
            in3 => \N__18672\,
            lcout => \QuadInstance3.Quad_RNO_0_2_1\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_0\,
            carryout => \QuadInstance3.un1_Quad_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_2_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30418\,
            in2 => \N__18828\,
            in3 => \N__18669\,
            lcout => \QuadInstance3.Quad_RNO_0_3_2\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_1\,
            carryout => \QuadInstance3.un1_Quad_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_3_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24367\,
            in2 => \N__18666\,
            in3 => \N__18654\,
            lcout => \QuadInstance3.Quad_RNO_0_3_3\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_2\,
            carryout => \QuadInstance3.un1_Quad_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_4_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19107\,
            in2 => \N__21845\,
            in3 => \N__18651\,
            lcout => \QuadInstance3.Quad_RNO_0_3_4\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_3\,
            carryout => \QuadInstance3.un1_Quad_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_5_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23741\,
            in2 => \N__18789\,
            in3 => \N__18777\,
            lcout => \QuadInstance3.Quad_RNO_0_3_5\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_4\,
            carryout => \QuadInstance3.un1_Quad_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_6_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28258\,
            in2 => \N__18774\,
            in3 => \N__18762\,
            lcout => \QuadInstance3.Quad_RNO_0_3_6\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_5\,
            carryout => \QuadInstance3.un1_Quad_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_7_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26329\,
            in2 => \N__19053\,
            in3 => \N__18759\,
            lcout => \QuadInstance3.Quad_RNO_0_3_7\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_6\,
            carryout => \QuadInstance3.un1_Quad_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_8_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30661\,
            in2 => \N__18807\,
            in3 => \N__18756\,
            lcout => \QuadInstance3.Quad_RNO_0_3_8\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \QuadInstance3.un1_Quad_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_9_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25480\,
            in2 => \N__18798\,
            in3 => \N__18753\,
            lcout => \QuadInstance3.Quad_RNO_0_3_9\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_8\,
            carryout => \QuadInstance3.un1_Quad_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_10_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34789\,
            in2 => \N__18816\,
            in3 => \N__18750\,
            lcout => \QuadInstance3.Quad_RNO_0_3_10\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_9\,
            carryout => \QuadInstance3.un1_Quad_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_11_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22414\,
            in2 => \N__18747\,
            in3 => \N__18738\,
            lcout => \QuadInstance3.Quad_RNO_0_3_11\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_10\,
            carryout => \QuadInstance3.un1_Quad_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_12_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22315\,
            in2 => \N__18735\,
            in3 => \N__18726\,
            lcout => \QuadInstance3.Quad_RNO_0_3_12\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_11\,
            carryout => \QuadInstance3.un1_Quad_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_13_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19928\,
            in2 => \N__18723\,
            in3 => \N__18714\,
            lcout => \QuadInstance3.Quad_RNO_0_3_13\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_12\,
            carryout => \QuadInstance3.un1_Quad_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_14_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19098\,
            in2 => \N__20072\,
            in3 => \N__18852\,
            lcout => \QuadInstance3.Quad_RNO_0_3_14\,
            ltout => OPEN,
            carryin => \QuadInstance3.un1_Quad_cry_13\,
            carryout => \QuadInstance3.un1_Quad_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_15_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__18888\,
            in1 => \N__21985\,
            in2 => \N__31908\,
            in3 => \N__18849\,
            lcout => \dataRead3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38609\,
            ce => 'H',
            sr => \N__35713\
        );

    \QuadInstance3.delayedCh_A_RNIO54L_2_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19074\,
            in1 => \N__19067\,
            in2 => \N__19089\,
            in3 => \N__18863\,
            lcout => \QuadInstance3.count_enable\,
            ltout => \QuadInstance3.count_enable_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNI8OAL1_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__23811\,
            in1 => \N__21917\,
            in2 => \N__18846\,
            in3 => \N__19022\,
            lcout => \QuadInstance3.Quad_RNI8OAL1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.delayedCh_B_RNIQUMH_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__34501\,
            in1 => \_gnd_net_\,
            in2 => \N__19088\,
            in3 => \N__19066\,
            lcout => \QuadInstance3.un1_count_enable_i_a2_0_1\,
            ltout => \QuadInstance3.un1_count_enable_i_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNI9PAL1_2_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__30422\,
            in1 => \N__21918\,
            in2 => \N__18831\,
            in3 => \N__18949\,
            lcout => \QuadInstance3.Quad_RNI9PAL1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIO10J1_10_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010110000"
        )
    port map (
            in0 => \N__21921\,
            in1 => \N__19034\,
            in2 => \N__18974\,
            in3 => \N__34803\,
            lcout => \QuadInstance3.Quad_RNIO10J1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIFVAL1_8_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__30668\,
            in1 => \N__21919\,
            in2 => \N__19040\,
            in3 => \N__18954\,
            lcout => \QuadInstance3.Quad_RNIFVAL1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIG0BL1_9_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010110000"
        )
    port map (
            in0 => \N__21920\,
            in1 => \N__19030\,
            in2 => \N__18973\,
            in3 => \N__25481\,
            lcout => \QuadInstance3.Quad_RNIG0BL1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIBRAL1_4_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001100"
        )
    port map (
            in0 => \N__21846\,
            in1 => \N__18950\,
            in2 => \N__21970\,
            in3 => \N__19023\,
            lcout => \QuadInstance3.Quad_RNIBRAL1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIS50J1_14_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__21934\,
            in1 => \N__18964\,
            in2 => \N__20079\,
            in3 => \N__19028\,
            lcout => \QuadInstance3.Quad_RNIS50J1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.delayedCh_B_2_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18864\,
            lcout => \QuadInstance3.delayedCh_BZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.delayedCh_A_2_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19068\,
            lcout => \QuadInstance3.delayedCh_AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.delayedCh_A_1_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20388\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance3.delayedCh_AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNIEUAL1_7_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__26336\,
            in1 => \N__21933\,
            in2 => \N__18975\,
            in3 => \N__19027\,
            lcout => \QuadInstance3.Quad_RNIEUAL1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.Quad_RNO_0_15_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010011100"
        )
    port map (
            in0 => \N__19029\,
            in1 => \N__24335\,
            in2 => \N__18977\,
            in3 => \N__21935\,
            lcout => \QuadInstance3.un1_Quad_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quadWrite_3_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__23444\,
            in1 => \N__33822\,
            in2 => \N__33661\,
            in3 => \N__33436\,
            lcout => \quadWriteZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance3.delayedCh_B_1_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18879\,
            lcout => \QuadInstance3.delayedCh_BZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__19179\,
            in1 => \N__19198\,
            in2 => \N__19394\,
            in3 => \N__19185\,
            lcout => \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.periodCounter_RNI5J7E_14_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__19255\,
            in1 => \N__19237\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \PWMInstance5.un1_periodCounter12_1_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.periodCounter_RNIIJIT_10_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19172\,
            in1 => \N__19219\,
            in2 => \N__19203\,
            in3 => \N__19199\,
            lcout => \PWMInstance5.un1_periodCounter12_1_0_a2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_4_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36494\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38578\,
            ce => \N__19597\,
            sr => \N__35739\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_5_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36366\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38578\,
            ce => \N__19597\,
            sr => \N__35739\
        );

    \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__19128\,
            in1 => \N__19171\,
            in2 => \N__19370\,
            in3 => \N__19158\,
            lcout => \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_11_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36004\,
            lcout => \PWMInstance5.PWMPulseWidthCountZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38578\,
            ce => \N__19597\,
            sr => \N__35739\
        );

    \PWMInstance5.out_RNO_0_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__19570\,
            in1 => \N__19552\,
            in2 => \N__20244\,
            in3 => \N__19316\,
            lcout => \PWMInstance5.un1_periodCounter12_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.clkCount_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100101"
        )
    port map (
            in0 => \N__19553\,
            in1 => \_gnd_net_\,
            in2 => \N__20231\,
            in3 => \N__19571\,
            lcout => \PWMInstance5.clkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38568\,
            ce => 'H',
            sr => \N__35747\
        );

    \PWMInstance5.PWMPulseWidthCount_esr_ctle_15_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35827\,
            in2 => \_gnd_net_\,
            in3 => \N__20224\,
            lcout => \PWMInstance5.pwmWrite_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.clkCount_1_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000001010"
        )
    port map (
            in0 => \N__19554\,
            in1 => \_gnd_net_\,
            in2 => \N__20232\,
            in3 => \N__19572\,
            lcout => \PWMInstance5.clkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38568\,
            ce => 'H',
            sr => \N__35747\
        );

    \PWMInstance5.clkCount_RNI8JO8_0_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__20240\,
            in1 => \N__19569\,
            in2 => \_gnd_net_\,
            in3 => \N__19551\,
            lcout => \PWMInstance5.periodCounter12\,
            ltout => \PWMInstance5.periodCounter12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.periodCounter_RNIP0851_15_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19519\,
            in1 => \N__19501\,
            in2 => \N__19482\,
            in3 => \N__19278\,
            lcout => OPEN,
            ltout => \PWMInstance5.un1_periodCounter12_1_0_a2_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.periodCounter_RNI8HQJ4_10_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19323\,
            in1 => \N__19479\,
            in2 => \N__19470\,
            in3 => \N__19467\,
            lcout => \PWMInstance5.out_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.periodCounter_RNIVUF81_11_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19414\,
            in1 => \N__19395\,
            in2 => \N__19371\,
            in3 => \N__19347\,
            lcout => \PWMInstance5.un1_periodCounter12_1_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance5.periodCounter_RNICQ7E_16_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19315\,
            in2 => \_gnd_net_\,
            in3 => \N__19299\,
            lcout => \PWMInstance5.un1_periodCounter12_1_0_a2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.periodCounter_RNI7M9F_14_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__23167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20210\,
            lcout => OPEN,
            ltout => \PWMInstance6.un1_periodCounter12_1_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.periodCounter_RNINBG41_10_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__23053\,
            in1 => \N__23128\,
            in2 => \N__19710\,
            in3 => \N__20351\,
            lcout => OPEN,
            ltout => \PWMInstance6.un1_periodCounter12_1_0_a2_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.periodCounter_RNISI7C4_10_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19704\,
            in1 => \N__21099\,
            in2 => \N__19707\,
            in3 => \N__21138\,
            lcout => \PWMInstance6.out_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.periodCounter_RNI34321_11_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21226\,
            in1 => \N__20323\,
            in2 => \N__23102\,
            in3 => \N__20179\,
            lcout => \PWMInstance6.un1_periodCounter12_1_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__19692\,
            in1 => \N__19698\,
            in2 => \N__20187\,
            in3 => \N__20211\,
            lcout => \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_2_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31592\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38550\,
            ce => \N__24556\,
            sr => \N__35763\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_3_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32072\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38550\,
            ce => \N__24556\,
            sr => \N__35763\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__20355\,
            in1 => \N__22959\,
            in2 => \N__19686\,
            in3 => \N__20328\,
            lcout => \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_4_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36512\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38550\,
            ce => \N__24556\,
            sr => \N__35763\
        );

    \QuadInstance2.Quad_2_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31587\,
            in1 => \N__22192\,
            in2 => \_gnd_net_\,
            in3 => \N__19677\,
            lcout => \dataRead2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38673\,
            ce => 'H',
            sr => \N__35690\
        );

    \QuadInstance3.Quad_2_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31589\,
            in1 => \N__22019\,
            in2 => \_gnd_net_\,
            in3 => \N__19665\,
            lcout => \dataRead3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38673\,
            ce => 'H',
            sr => \N__35690\
        );

    \QuadInstance2.Quad_6_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31120\,
            in1 => \N__22194\,
            in2 => \_gnd_net_\,
            in3 => \N__19770\,
            lcout => \dataRead2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38673\,
            ce => 'H',
            sr => \N__35690\
        );

    \QuadInstance6.Quad_2_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31590\,
            in1 => \N__22798\,
            in2 => \_gnd_net_\,
            in3 => \N__20430\,
            lcout => \dataRead6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38673\,
            ce => 'H',
            sr => \N__35690\
        );

    \QuadInstance7.Quad_2_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31588\,
            in1 => \N__26052\,
            in2 => \_gnd_net_\,
            in3 => \N__19758\,
            lcout => \dataRead7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38673\,
            ce => 'H',
            sr => \N__35690\
        );

    \QuadInstance1.Quad_3_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24098\,
            in1 => \N__32086\,
            in2 => \_gnd_net_\,
            in3 => \N__21615\,
            lcout => \dataRead1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38673\,
            ce => 'H',
            sr => \N__35690\
        );

    \QuadInstance2.Quad_3_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32087\,
            in1 => \N__22193\,
            in2 => \_gnd_net_\,
            in3 => \N__19746\,
            lcout => \dataRead2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38673\,
            ce => 'H',
            sr => \N__35690\
        );

    \QuadInstance5.Quad_4_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36514\,
            in1 => \N__25800\,
            in2 => \_gnd_net_\,
            in3 => \N__19734\,
            lcout => \dataRead5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38662\,
            ce => 'H',
            sr => \N__35692\
        );

    \QuadInstance5.Quad_6_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25798\,
            in1 => \N__31112\,
            in2 => \_gnd_net_\,
            in3 => \N__19728\,
            lcout => \dataRead5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38662\,
            ce => 'H',
            sr => \N__35692\
        );

    \QuadInstance6.Quad_6_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31113\,
            in1 => \N__22796\,
            in2 => \_gnd_net_\,
            in3 => \N__20508\,
            lcout => \dataRead6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38662\,
            ce => 'H',
            sr => \N__35692\
        );

    \QuadInstance7.Quad_6_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31110\,
            in1 => \N__26014\,
            in2 => \_gnd_net_\,
            in3 => \N__19722\,
            lcout => \dataRead7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38662\,
            ce => 'H',
            sr => \N__35692\
        );

    \QuadInstance7.Quad_9_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26013\,
            in1 => \N__28572\,
            in2 => \_gnd_net_\,
            in3 => \N__19836\,
            lcout => \dataRead7_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38662\,
            ce => 'H',
            sr => \N__35692\
        );

    \QuadInstance5.Quad_8_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25799\,
            in1 => \N__28988\,
            in2 => \_gnd_net_\,
            in3 => \N__19824\,
            lcout => \dataRead5_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38662\,
            ce => 'H',
            sr => \N__35692\
        );

    \QuadInstance6.Quad_8_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28989\,
            in1 => \N__22797\,
            in2 => \_gnd_net_\,
            in3 => \N__20490\,
            lcout => \dataRead6_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38662\,
            ce => 'H',
            sr => \N__35692\
        );

    \QuadInstance3.Quad_3_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32073\,
            in1 => \N__22018\,
            in2 => \_gnd_net_\,
            in3 => \N__19815\,
            lcout => \dataRead3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38662\,
            ce => 'H',
            sr => \N__35692\
        );

    \QuadInstance1.Quad_7_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29448\,
            in1 => \_gnd_net_\,
            in2 => \N__24099\,
            in3 => \N__21564\,
            lcout => \dataRead1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38650\,
            ce => 'H',
            sr => \N__35700\
        );

    \QuadInstance2.Quad_7_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29449\,
            in1 => \N__22185\,
            in2 => \_gnd_net_\,
            in3 => \N__19803\,
            lcout => \dataRead2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38650\,
            ce => 'H',
            sr => \N__35700\
        );

    \QuadInstance3.Quad_7_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22015\,
            in1 => \N__29450\,
            in2 => \_gnd_net_\,
            in3 => \N__19794\,
            lcout => \dataRead3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38650\,
            ce => 'H',
            sr => \N__35700\
        );

    \QuadInstance5.Quad_7_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29451\,
            in1 => \N__25772\,
            in2 => \_gnd_net_\,
            in3 => \N__19785\,
            lcout => \dataRead5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38650\,
            ce => 'H',
            sr => \N__35700\
        );

    \QuadInstance3.Quad_5_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22014\,
            in1 => \N__36368\,
            in2 => \_gnd_net_\,
            in3 => \N__19779\,
            lcout => \dataRead3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38650\,
            ce => 'H',
            sr => \N__35700\
        );

    \QuadInstance7.Quad_7_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29452\,
            in1 => \N__26012\,
            in2 => \_gnd_net_\,
            in3 => \N__19890\,
            lcout => \dataRead7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38650\,
            ce => 'H',
            sr => \N__35700\
        );

    \QuadInstance1.Quad_8_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24080\,
            in1 => \N__28987\,
            in2 => \_gnd_net_\,
            in3 => \N__21552\,
            lcout => \dataRead1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38650\,
            ce => 'H',
            sr => \N__35700\
        );

    \QuadInstance6.Quad_11_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__35993\,
            in1 => \_gnd_net_\,
            in2 => \N__22805\,
            in3 => \N__20475\,
            lcout => \dataRead6_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38650\,
            ce => 'H',
            sr => \N__35700\
        );

    \QuadInstance0.Quad_11_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36005\,
            in1 => \N__33132\,
            in2 => \_gnd_net_\,
            in3 => \N__30066\,
            lcout => \dataRead0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38641\,
            ce => 'H',
            sr => \N__35705\
        );

    \QuadInstance1.Quad_11_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24095\,
            in1 => \N__36006\,
            in2 => \_gnd_net_\,
            in3 => \N__21675\,
            lcout => \dataRead1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38641\,
            ce => 'H',
            sr => \N__35705\
        );

    \QuadInstance2.Quad_11_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22186\,
            in1 => \_gnd_net_\,
            in2 => \N__36015\,
            in3 => \N__19878\,
            lcout => \dataRead2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38641\,
            ce => 'H',
            sr => \N__35705\
        );

    \QuadInstance5.Quad_10_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25796\,
            in1 => \N__36142\,
            in2 => \_gnd_net_\,
            in3 => \N__19869\,
            lcout => \dataRead5_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38641\,
            ce => 'H',
            sr => \N__35705\
        );

    \QuadInstance5.Quad_11_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36010\,
            in1 => \N__25797\,
            in2 => \_gnd_net_\,
            in3 => \N__19863\,
            lcout => \dataRead5_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38641\,
            ce => 'H',
            sr => \N__35705\
        );

    \QuadInstance2.Quad_8_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28986\,
            in1 => \N__22187\,
            in2 => \_gnd_net_\,
            in3 => \N__19857\,
            lcout => \dataRead2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38641\,
            ce => 'H',
            sr => \N__35705\
        );

    \QuadInstance3.Quad_9_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28559\,
            in1 => \N__22017\,
            in2 => \_gnd_net_\,
            in3 => \N__19845\,
            lcout => \dataRead3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38641\,
            ce => 'H',
            sr => \N__35705\
        );

    \QuadInstance0.Quad_3_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33131\,
            in1 => \N__32050\,
            in2 => \_gnd_net_\,
            in3 => \N__29865\,
            lcout => \dataRead0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38641\,
            ce => 'H',
            sr => \N__35705\
        );

    \OutReg_ess_RNO_3_13_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__28013\,
            in1 => \N__19921\,
            in2 => \N__28133\,
            in3 => \N__19960\,
            lcout => \OutReg_0_4_i_m3_ns_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_2_13_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__23922\,
            in1 => \N__38152\,
            in2 => \N__20019\,
            in3 => \N__27543\,
            lcout => \OutReg_ess_RNO_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.Quad_13_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28684\,
            in1 => \N__22188\,
            in2 => \_gnd_net_\,
            in3 => \N__19986\,
            lcout => \dataRead2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38631\,
            ce => 'H',
            sr => \N__35714\
        );

    \QuadInstance3.Quad_13_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22016\,
            in1 => \N__28685\,
            in2 => \_gnd_net_\,
            in3 => \N__19944\,
            lcout => \dataRead3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38631\,
            ce => 'H',
            sr => \N__35714\
        );

    \QuadInstance6.Quad_13_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28686\,
            in1 => \N__22755\,
            in2 => \_gnd_net_\,
            in3 => \N__20625\,
            lcout => \dataRead6_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38631\,
            ce => 'H',
            sr => \N__35714\
        );

    \QuadInstance3.Quad_12_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28800\,
            in1 => \N__22003\,
            in2 => \_gnd_net_\,
            in3 => \N__19905\,
            lcout => \dataRead3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38618\,
            ce => 'H',
            sr => \N__35721\
        );

    \QuadInstance6.Quad_12_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28801\,
            in1 => \N__22754\,
            in2 => \_gnd_net_\,
            in3 => \N__20466\,
            lcout => \dataRead6_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38618\,
            ce => 'H',
            sr => \N__35721\
        );

    \QuadInstance3.Quad_8_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28952\,
            in1 => \_gnd_net_\,
            in2 => \N__19899\,
            in3 => \N__22004\,
            lcout => \dataRead3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38618\,
            ce => 'H',
            sr => \N__35721\
        );

    \QuadInstance3.Quad_14_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22000\,
            in1 => \N__34365\,
            in2 => \_gnd_net_\,
            in3 => \N__20157\,
            lcout => \dataRead3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38618\,
            ce => 'H',
            sr => \N__35721\
        );

    \QuadInstance5.Quad_2_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31542\,
            in1 => \N__25806\,
            in2 => \_gnd_net_\,
            in3 => \N__20151\,
            lcout => \dataRead5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38618\,
            ce => 'H',
            sr => \N__35721\
        );

    \QuadInstance7.Quad_14_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34366\,
            in1 => \N__26038\,
            in2 => \_gnd_net_\,
            in3 => \N__20142\,
            lcout => \dataRead7_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38618\,
            ce => 'H',
            sr => \N__35721\
        );

    \QuadInstance3.Quad_10_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36089\,
            in1 => \N__22002\,
            in2 => \_gnd_net_\,
            in3 => \N__20133\,
            lcout => \dataRead3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38618\,
            ce => 'H',
            sr => \N__35721\
        );

    \QuadInstance3.Quad_11_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22001\,
            in1 => \_gnd_net_\,
            in2 => \N__35973\,
            in3 => \N__20127\,
            lcout => \dataRead3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38618\,
            ce => 'H',
            sr => \N__35721\
        );

    \OutReg_ess_RNO_0_13_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37558\,
            in1 => \N__20121\,
            in2 => \_gnd_net_\,
            in3 => \N__20730\,
            lcout => \OutReg_ess_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_4_11_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__28015\,
            in1 => \N__30097\,
            in2 => \N__25122\,
            in3 => \N__28137\,
            lcout => OPEN,
            ltout => \OutReg_0_5_i_m3_i_m3_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_2_11_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__20108\,
            in1 => \N__32948\,
            in2 => \N__20082\,
            in3 => \N__23366\,
            lcout => \OutReg_ess_RNO_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_3_14_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__20065\,
            in1 => \N__20048\,
            in2 => \N__28140\,
            in3 => \N__28014\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_1_14_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__20263\,
            in1 => \N__20558\,
            in2 => \N__20247\,
            in3 => \N__37741\,
            lcout => \OutReg_esr_RNO_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33749\,
            in1 => \N__33560\,
            in2 => \N__33464\,
            in3 => \N__33207\,
            lcout => \pwmWriteZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_esr_4_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30621\,
            lcout => \data_receivedZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38590\,
            ce => \N__26184\,
            sr => \N__26154\
        );

    \pwmWrite_fast_5_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__23429\,
            in1 => \N__33440\,
            in2 => \N__33600\,
            in3 => \N__33751\,
            lcout => \pwmWrite_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_5_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33750\,
            in1 => \N__33561\,
            in2 => \N__33465\,
            in3 => \N__23428\,
            lcout => \pwmWriteZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.periodCounter_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21090\,
            in2 => \N__21162\,
            in3 => \N__21158\,
            lcout => \PWMInstance6.periodCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_0\,
            clk => \N__38569\,
            ce => 'H',
            sr => \N__35298\
        );

    \PWMInstance6.periodCounter_1_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21074\,
            in2 => \_gnd_net_\,
            in3 => \N__20214\,
            lcout => \PWMInstance6.periodCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_0\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_1\,
            clk => \N__38569\,
            ce => 'H',
            sr => \N__35298\
        );

    \PWMInstance6.periodCounter_2_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20209\,
            in2 => \_gnd_net_\,
            in3 => \N__20190\,
            lcout => \PWMInstance6.periodCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_1\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_2\,
            clk => \N__38569\,
            ce => 'H',
            sr => \N__35298\
        );

    \PWMInstance6.periodCounter_3_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20180\,
            in2 => \_gnd_net_\,
            in3 => \N__20160\,
            lcout => \PWMInstance6.periodCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_2\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_3\,
            clk => \N__38569\,
            ce => 'H',
            sr => \N__35298\
        );

    \PWMInstance6.periodCounter_4_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20350\,
            in2 => \_gnd_net_\,
            in3 => \N__20331\,
            lcout => \PWMInstance6.periodCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_3\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_4\,
            clk => \N__38569\,
            ce => 'H',
            sr => \N__35298\
        );

    \PWMInstance6.periodCounter_5_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20327\,
            in2 => \_gnd_net_\,
            in3 => \N__20307\,
            lcout => \PWMInstance6.periodCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_4\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_5\,
            clk => \N__38569\,
            ce => 'H',
            sr => \N__35298\
        );

    \PWMInstance6.periodCounter_6_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21041\,
            in2 => \_gnd_net_\,
            in3 => \N__20304\,
            lcout => \PWMInstance6.periodCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_5\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_6\,
            clk => \N__38569\,
            ce => 'H',
            sr => \N__35298\
        );

    \PWMInstance6.periodCounter_7_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21422\,
            in1 => \N__21024\,
            in2 => \_gnd_net_\,
            in3 => \N__20301\,
            lcout => \PWMInstance6.periodCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_6\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_7\,
            clk => \N__38569\,
            ce => 'H',
            sr => \N__35298\
        );

    \PWMInstance6.periodCounter_8_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21246\,
            in2 => \_gnd_net_\,
            in3 => \N__20298\,
            lcout => \PWMInstance6.periodCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_8\,
            clk => \N__38562\,
            ce => 'H',
            sr => \N__35296\
        );

    \PWMInstance6.periodCounter_9_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21227\,
            in2 => \_gnd_net_\,
            in3 => \N__20295\,
            lcout => \PWMInstance6.periodCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_8\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_9\,
            clk => \N__38562\,
            ce => 'H',
            sr => \N__35296\
        );

    \PWMInstance6.periodCounter_10_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23129\,
            in2 => \_gnd_net_\,
            in3 => \N__20292\,
            lcout => \PWMInstance6.periodCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_9\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_10\,
            clk => \N__38562\,
            ce => 'H',
            sr => \N__35296\
        );

    \PWMInstance6.periodCounter_11_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21420\,
            in1 => \N__23098\,
            in2 => \_gnd_net_\,
            in3 => \N__20289\,
            lcout => \PWMInstance6.periodCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_10\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_11\,
            clk => \N__38562\,
            ce => 'H',
            sr => \N__35296\
        );

    \PWMInstance6.periodCounter_12_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21412\,
            in1 => \N__23054\,
            in2 => \_gnd_net_\,
            in3 => \N__20286\,
            lcout => \PWMInstance6.periodCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_11\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_12\,
            clk => \N__38562\,
            ce => 'H',
            sr => \N__35296\
        );

    \PWMInstance6.periodCounter_13_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21421\,
            in1 => \N__23030\,
            in2 => \_gnd_net_\,
            in3 => \N__20412\,
            lcout => \PWMInstance6.periodCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_12\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_13\,
            clk => \N__38562\,
            ce => 'H',
            sr => \N__35296\
        );

    \PWMInstance6.periodCounter_14_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23175\,
            in2 => \_gnd_net_\,
            in3 => \N__20409\,
            lcout => \PWMInstance6.periodCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_13\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_14\,
            clk => \N__38562\,
            ce => 'H',
            sr => \N__35296\
        );

    \PWMInstance6.periodCounter_15_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23196\,
            in2 => \_gnd_net_\,
            in3 => \N__20406\,
            lcout => \PWMInstance6.periodCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_periodCounter_2_cry_14\,
            carryout => \PWMInstance6.un1_periodCounter_2_cry_15\,
            clk => \N__38562\,
            ce => 'H',
            sr => \N__35296\
        );

    \PWMInstance6.periodCounter_16_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21413\,
            in1 => \N__20923\,
            in2 => \_gnd_net_\,
            in3 => \N__20403\,
            lcout => \PWMInstance6.periodCounterZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38555\,
            ce => 'H',
            sr => \N__35294\
        );

    \QuadInstance3.delayedCh_A_0_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20400\,
            lcout => \QuadInstance3.delayedCh_AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38702\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNIKINB1_14_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__22791\,
            in1 => \N__22634\,
            in2 => \N__20562\,
            in3 => \N__22562\,
            lcout => \QuadInstance6.Quad_RNIKINB1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_15_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111110000"
        )
    port map (
            in0 => \N__22792\,
            in1 => \N__22635\,
            in2 => \N__24273\,
            in3 => \N__22563\,
            lcout => \QuadInstance6.un1_Quad_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_5_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__24100\,
            in1 => \N__21591\,
            in2 => \_gnd_net_\,
            in3 => \N__36371\,
            lcout => \dataRead1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38680\,
            ce => 'H',
            sr => \N__35693\
        );

    \QuadInstance2.Quad_5_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22191\,
            in1 => \_gnd_net_\,
            in2 => \N__36378\,
            in3 => \N__20370\,
            lcout => \dataRead2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38680\,
            ce => 'H',
            sr => \N__35693\
        );

    \QuadInstance6.Quad_7_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22794\,
            in1 => \_gnd_net_\,
            in2 => \N__29443\,
            in3 => \N__20499\,
            lcout => \dataRead6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38680\,
            ce => 'H',
            sr => \N__35693\
        );

    \QuadInstance5.Quad_5_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36369\,
            in1 => \N__25795\,
            in2 => \_gnd_net_\,
            in3 => \N__20457\,
            lcout => \dataRead5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38680\,
            ce => 'H',
            sr => \N__35693\
        );

    \QuadInstance6.Quad_5_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22793\,
            in1 => \N__36372\,
            in2 => \_gnd_net_\,
            in3 => \N__20517\,
            lcout => \dataRead6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38680\,
            ce => 'H',
            sr => \N__35693\
        );

    \QuadInstance7.Quad_5_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36370\,
            in1 => \N__26053\,
            in2 => \_gnd_net_\,
            in3 => \N__20445\,
            lcout => \dataRead7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38680\,
            ce => 'H',
            sr => \N__35693\
        );

    \QuadInstance1.Quad_6_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__24101\,
            in1 => \N__31111\,
            in2 => \N__21579\,
            in3 => \_gnd_net_\,
            lcout => \dataRead1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38680\,
            ce => 'H',
            sr => \N__35693\
        );

    \QuadInstance6.Quad_3_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32083\,
            in1 => \N__22795\,
            in2 => \_gnd_net_\,
            in3 => \N__20421\,
            lcout => \dataRead6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38680\,
            ce => 'H',
            sr => \N__35693\
        );

    \QuadInstance6.un1_Quad_cry_0_c_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22555\,
            in2 => \N__30810\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \QuadInstance6.un1_Quad_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_1_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23783\,
            in2 => \N__20703\,
            in3 => \N__20433\,
            lcout => \QuadInstance6.Quad_RNO_0_5_1\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_0\,
            carryout => \QuadInstance6.un1_Quad_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_2_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30346\,
            in2 => \N__20688\,
            in3 => \N__20424\,
            lcout => \QuadInstance6.Quad_RNO_0_6_2\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_1\,
            carryout => \QuadInstance6.un1_Quad_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_3_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27796\,
            in2 => \N__20664\,
            in3 => \N__20415\,
            lcout => \QuadInstance6.Quad_RNO_0_6_3\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_2\,
            carryout => \QuadInstance6.un1_Quad_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21500\,
            in2 => \N__20784\,
            in3 => \N__20520\,
            lcout => \QuadInstance6.Quad_RNO_0_6_4\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_3\,
            carryout => \QuadInstance6.un1_Quad_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_5_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36766\,
            in2 => \N__20652\,
            in3 => \N__20511\,
            lcout => \QuadInstance6.Quad_RNO_0_6_5\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_4\,
            carryout => \QuadInstance6.un1_Quad_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27724\,
            in2 => \N__20760\,
            in3 => \N__20502\,
            lcout => \QuadInstance6.Quad_RNO_0_6_6\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_5\,
            carryout => \QuadInstance6.un1_Quad_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_7_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26287\,
            in2 => \N__20748\,
            in3 => \N__20493\,
            lcout => \QuadInstance6.Quad_RNO_0_6_7\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_6\,
            carryout => \QuadInstance6.un1_Quad_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_8_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37783\,
            in2 => \N__20799\,
            in3 => \N__20484\,
            lcout => \QuadInstance6.Quad_RNO_0_6_8\,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \QuadInstance6.un1_Quad_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_9_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25419\,
            in2 => \N__20640\,
            in3 => \N__20481\,
            lcout => \QuadInstance6.Quad_RNO_0_6_9\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_8\,
            carryout => \QuadInstance6.un1_Quad_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_10_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34609\,
            in2 => \N__21702\,
            in3 => \N__20478\,
            lcout => \QuadInstance6.Quad_RNO_0_6_10\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_9\,
            carryout => \QuadInstance6.un1_Quad_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_11_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20830\,
            in2 => \N__20676\,
            in3 => \N__20469\,
            lcout => \QuadInstance6.Quad_RNO_0_6_11\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_10\,
            carryout => \QuadInstance6.un1_Quad_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_12_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22289\,
            in2 => \N__20772\,
            in3 => \N__20628\,
            lcout => \QuadInstance6.Quad_RNO_0_6_12\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_11\,
            carryout => \QuadInstance6.un1_Quad_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_13_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22476\,
            in2 => \N__22839\,
            in3 => \N__20616\,
            lcout => \QuadInstance6.Quad_RNO_0_6_13\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_12\,
            carryout => \QuadInstance6.un1_Quad_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNO_0_14_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20613\,
            in2 => \N__20554\,
            in3 => \N__20604\,
            lcout => \QuadInstance6.Quad_RNO_0_6_14\,
            ltout => OPEN,
            carryin => \QuadInstance6.un1_Quad_cry_13\,
            carryout => \QuadInstance6.un1_Quad_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_15_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__22783\,
            in1 => \N__20601\,
            in2 => \N__31895\,
            in3 => \N__20592\,
            lcout => \dataRead6_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38663\,
            ce => 'H',
            sr => \N__35706\
        );

    \QuadInstance1.Quad_10_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36133\,
            in1 => \N__24096\,
            in2 => \_gnd_net_\,
            in3 => \N__21684\,
            lcout => \dataRead1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38651\,
            ce => 'H',
            sr => \N__35715\
        );

    \QuadInstance6.Quad_1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22788\,
            in1 => \N__31247\,
            in2 => \_gnd_net_\,
            in3 => \N__20589\,
            lcout => \dataRead6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38651\,
            ce => 'H',
            sr => \N__35715\
        );

    \QuadInstance7.Quad_8_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26054\,
            in1 => \N__28985\,
            in2 => \_gnd_net_\,
            in3 => \N__20580\,
            lcout => \dataRead7_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38651\,
            ce => 'H',
            sr => \N__35715\
        );

    \QuadInstance6.Quad_14_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22787\,
            in1 => \N__34374\,
            in2 => \_gnd_net_\,
            in3 => \N__20568\,
            lcout => \dataRead6_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38651\,
            ce => 'H',
            sr => \N__35715\
        );

    \QuadInstance6.Quad_10_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36134\,
            in1 => \N__22789\,
            in2 => \_gnd_net_\,
            in3 => \N__20526\,
            lcout => \dataRead6_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38651\,
            ce => 'H',
            sr => \N__35715\
        );

    \QuadInstance7.Quad_10_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36135\,
            in1 => \N__26055\,
            in2 => \_gnd_net_\,
            in3 => \N__20724\,
            lcout => \dataRead7_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38651\,
            ce => 'H',
            sr => \N__35715\
        );

    \QuadInstance1.Quad_14_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34373\,
            in1 => \N__24097\,
            in2 => \_gnd_net_\,
            in3 => \N__21657\,
            lcout => \dataRead1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38651\,
            ce => 'H',
            sr => \N__35715\
        );

    \QuadInstance5.Quad_9_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28558\,
            in1 => \N__25802\,
            in2 => \_gnd_net_\,
            in3 => \N__20712\,
            lcout => \dataRead5_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38651\,
            ce => 'H',
            sr => \N__35715\
        );

    \QuadInstance6.Quad_RNI02A91_1_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__23782\,
            in1 => \N__22704\,
            in2 => \N__22551\,
            in3 => \N__22604\,
            lcout => \QuadInstance6.Quad_RNI02A91Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.delayedCh_A_RNI4QLG_2_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22466\,
            in1 => \N__22862\,
            in2 => \N__21720\,
            in3 => \N__22845\,
            lcout => \QuadInstance6.count_enable\,
            ltout => \QuadInstance6.count_enable_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNI13A91_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__30354\,
            in1 => \N__22705\,
            in2 => \N__20691\,
            in3 => \N__22605\,
            lcout => \QuadInstance6.Quad_RNI13A91Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNIHFNB1_11_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000100"
        )
    port map (
            in0 => \N__22610\,
            in1 => \N__22533\,
            in2 => \N__22758\,
            in3 => \N__20840\,
            lcout => \QuadInstance6.Quad_RNIHFNB1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNI24A91_3_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__27812\,
            in1 => \N__22706\,
            in2 => \N__22552\,
            in3 => \N__22606\,
            lcout => \QuadInstance6.Quad_RNI24A91Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNI46A91_5_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__22607\,
            in1 => \N__36776\,
            in2 => \N__22756\,
            in3 => \N__22528\,
            lcout => \QuadInstance6.Quad_RNI46A91Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNI8AA91_9_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__25418\,
            in1 => \N__22710\,
            in2 => \N__22553\,
            in3 => \N__22609\,
            lcout => \QuadInstance6.Quad_RNI8AA91Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNI79A91_8_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__22608\,
            in1 => \N__37787\,
            in2 => \N__22757\,
            in3 => \N__22529\,
            lcout => \QuadInstance6.Quad_RNI79A91Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.delayedCh_B_RNI0PFF_2_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34469\,
            in2 => \N__21719\,
            in3 => \N__22861\,
            lcout => \QuadInstance6.un1_count_enable_i_a2_0_1\,
            ltout => \QuadInstance6.un1_count_enable_i_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNI35A91_4_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__21504\,
            in1 => \N__22717\,
            in2 => \N__20787\,
            in3 => \N__22534\,
            lcout => \QuadInstance6.Quad_RNI35A91Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.delayedCh_A_1_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21111\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance6.delayedCh_AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38632\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNIIGNB1_12_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__22282\,
            in1 => \N__22720\,
            in2 => \N__22631\,
            in3 => \N__22539\,
            lcout => \QuadInstance6.Quad_RNIIGNB1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNI57A91_6_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__22719\,
            in1 => \N__27740\,
            in2 => \N__22554\,
            in3 => \N__22614\,
            lcout => \QuadInstance6.Quad_RNI57A91Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNI68A91_7_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__26303\,
            in1 => \N__22718\,
            in2 => \N__22630\,
            in3 => \N__22538\,
            lcout => \QuadInstance6.Quad_RNI68A91Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_13_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010101"
        )
    port map (
            in0 => \N__20736\,
            in1 => \N__22822\,
            in2 => \N__26107\,
            in3 => \N__37748\,
            lcout => \OutReg_ess_RNO_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quadWrite_6_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33826\,
            in1 => \N__33599\,
            in2 => \N__33467\,
            in3 => \N__33203\,
            lcout => \quadWriteZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38632\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_11_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001010101"
        )
    port map (
            in0 => \N__22395\,
            in1 => \N__20876\,
            in2 => \N__20844\,
            in3 => \N__32839\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_1Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_0_11_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37560\,
            in2 => \N__20817\,
            in3 => \N__20814\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_0Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_11_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__34911\,
            in1 => \N__38883\,
            in2 => \N__20808\,
            in3 => \N__37394\,
            lcout => \OutRegZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38619\,
            ce => \N__37251\,
            sr => \N__37133\
        );

    \OutReg_ess_13_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__37395\,
            in1 => \N__20805\,
            in2 => \N__38911\,
            in3 => \N__22929\,
            lcout => \OutRegZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38619\,
            ce => \N__37251\,
            sr => \N__37133\
        );

    \dataWrite_0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38157\,
            lcout => \dataWriteZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \dataWrite_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37563\,
            lcout => \dataWriteZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \dataWrite_10_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22887\,
            lcout => \dataWriteZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \dataWrite_11_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22875\,
            lcout => \dataWriteZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \dataWrite_12_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22923\,
            lcout => \dataWriteZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \dataWrite_13_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22911\,
            lcout => \dataWriteZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \dataWrite_14_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22898\,
            lcout => \dataWriteZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \dataWrite_15_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20889\,
            lcout => \dataWriteZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__24461\,
            sr => \_gnd_net_\
        );

    \data_received_esr_18_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20901\,
            lcout => \data_receivedZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38598\,
            ce => \N__26181\,
            sr => \N__26151\
        );

    \data_received_esr_19_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20907\,
            lcout => \data_receivedZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38598\,
            ce => \N__26181\,
            sr => \N__26151\
        );

    \data_received_esr_20_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22995\,
            lcout => \data_receivedZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38598\,
            ce => \N__26181\,
            sr => \N__26151\
        );

    \data_received_esr_17_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20895\,
            lcout => \data_receivedZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38598\,
            ce => \N__26181\,
            sr => \N__26151\
        );

    \data_received_esr_16_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20888\,
            lcout => \data_receivedZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38598\,
            ce => \N__26181\,
            sr => \N__26151\
        );

    \data_received_esr_15_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22899\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \data_receivedZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38598\,
            ce => \N__26181\,
            sr => \N__26151\
        );

    \data_received_esr_3_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37764\,
            lcout => \data_receivedZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38598\,
            ce => \N__26181\,
            sr => \N__26151\
        );

    \data_received_esr_21_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33586\,
            lcout => \data_receivedZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38598\,
            ce => \N__26181\,
            sr => \N__26151\
        );

    \PWMInstance6.clkCount_0_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__20942\,
            in1 => \N__20969\,
            in2 => \_gnd_net_\,
            in3 => \N__20990\,
            lcout => \PWMInstance6.clkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38591\,
            ce => 'H',
            sr => \N__35757\
        );

    \PWMInstance6.clkCount_1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001011000010"
        )
    port map (
            in0 => \N__20991\,
            in1 => \N__20943\,
            in2 => \N__20973\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance6.clkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38591\,
            ce => 'H',
            sr => \N__35757\
        );

    \PWMInstance6.out_RNO_0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20952\,
            in1 => \N__20989\,
            in2 => \N__20928\,
            in3 => \N__20968\,
            lcout => \PWMInstance6.un1_periodCounter12_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_6_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33192\,
            in1 => \N__33456\,
            in2 => \N__33637\,
            in3 => \N__33783\,
            lcout => \pwmWriteZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.clkCount_RNIBCT4_0_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__20951\,
            in1 => \N__20988\,
            in2 => \_gnd_net_\,
            in3 => \N__20967\,
            lcout => \PWMInstance6.periodCounter12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_fast_6_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33193\,
            in1 => \N__33457\,
            in2 => \N__33638\,
            in3 => \N__33784\,
            lcout => \pwmWrite_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_ctle_15_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__35829\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20941\,
            lcout => \PWMInstance6.pwmWrite_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.periodCounter_RNIET9F_16_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20924\,
            in2 => \_gnd_net_\,
            in3 => \N__21022\,
            lcout => OPEN,
            ltout => \PWMInstance6.un1_periodCounter12_1_0_a2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.periodCounter_RNI00H31_15_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21073\,
            in1 => \N__23188\,
            in2 => \N__21165\,
            in3 => \N__21154\,
            lcout => \PWMInstance6.un1_periodCounter12_1_0_a2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.delayedCh_A_0_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21126\,
            lcout => \QuadInstance6.delayedCh_AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.periodCounter_RNI23321_13_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21089\,
            in1 => \N__23026\,
            in2 => \N__21042\,
            in3 => \N__21245\,
            lcout => \PWMInstance6.un1_periodCounter12_1_0_a2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__21048\,
            in1 => \N__21088\,
            in2 => \N__21075\,
            in3 => \N__21054\,
            lcout => \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_0_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31378\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38570\,
            ce => \N__24557\,
            sr => \N__35769\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_1_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31257\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38570\,
            ce => \N__24557\,
            sr => \N__35769\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__21037\,
            in1 => \N__21006\,
            in2 => \N__21000\,
            in3 => \N__21023\,
            lcout => \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_6_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31119\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38570\,
            ce => \N__24557\,
            sr => \N__35769\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_7_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29444\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38570\,
            ce => \N__24557\,
            sr => \N__35769\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__22947\,
            in1 => \N__21244\,
            in2 => \N__21228\,
            in3 => \N__24570\,
            lcout => \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21207\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32314\,
            in2 => \N__21201\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_0\,
            carryout => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21189\,
            in2 => \N__32410\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_1\,
            carryout => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32306\,
            in2 => \N__21180\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_2\,
            carryout => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21171\,
            in2 => \N__32412\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_3\,
            carryout => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32307\,
            in2 => \N__23076\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_4\,
            carryout => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23004\,
            in2 => \N__32411\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_5\,
            carryout => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32305\,
            in2 => \N__23154\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_6\,
            carryout => \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.out_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__21368\,
            in1 => \N__21435\,
            in2 => \N__21426\,
            in3 => \N__21381\,
            lcout => \PWM6_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38556\,
            ce => 'H',
            sr => \N__35781\
        );

    \PWM5_obufLegalizeSB_DFF_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM5_obufLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance2.delayedCh_A_0_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21351\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance2.delayedCh_AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_1_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24059\,
            in1 => \N__31271\,
            in2 => \_gnd_net_\,
            in3 => \N__21645\,
            lcout => \dataRead1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38695\,
            ce => 'H',
            sr => \N__35694\
        );

    \OutReg_ess_RNO_2_4_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__21327\,
            in1 => \N__38153\,
            in2 => \N__23265\,
            in3 => \N__21252\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_0_4_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37556\,
            in2 => \N__21300\,
            in3 => \N__21258\,
            lcout => \OutReg_ess_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_3_4_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__34763\,
            in1 => \N__21838\,
            in2 => \N__34896\,
            in3 => \N__21295\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_4_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__21496\,
            in1 => \N__21451\,
            in2 => \N__21261\,
            in3 => \N__37737\,
            lcout => \OutReg_ess_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_4_4_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__34153\,
            in1 => \N__28138\,
            in2 => \N__28017\,
            in3 => \N__27517\,
            lcout => \OutReg_0_5_i_m3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.delayedCh_A_0_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21540\,
            lcout => \QuadInstance0.delayedCh_AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_4_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33128\,
            in1 => \N__36484\,
            in2 => \_gnd_net_\,
            in3 => \N__29847\,
            lcout => \dataRead0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38681\,
            ce => 'H',
            sr => \N__35707\
        );

    \QuadInstance1.Quad_4_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36485\,
            in1 => \N__24051\,
            in2 => \_gnd_net_\,
            in3 => \N__21600\,
            lcout => \dataRead1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38681\,
            ce => 'H',
            sr => \N__35707\
        );

    \QuadInstance4.Quad_1_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29658\,
            in1 => \N__31252\,
            in2 => \_gnd_net_\,
            in3 => \N__24951\,
            lcout => \dataRead4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38681\,
            ce => 'H',
            sr => \N__35707\
        );

    \QuadInstance4.Quad_4_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36486\,
            in1 => \N__29659\,
            in2 => \_gnd_net_\,
            in3 => \N__24930\,
            lcout => \dataRead4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38681\,
            ce => 'H',
            sr => \N__35707\
        );

    \QuadInstance3.Quad_6_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31109\,
            in1 => \N__22020\,
            in2 => \_gnd_net_\,
            in3 => \N__21525\,
            lcout => \dataRead3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38681\,
            ce => 'H',
            sr => \N__35707\
        );

    \QuadInstance6.Quad_4_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__36487\,
            in1 => \N__22806\,
            in2 => \N__21513\,
            in3 => \_gnd_net_\,
            lcout => \dataRead6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38681\,
            ce => 'H',
            sr => \N__35707\
        );

    \QuadInstance7.Quad_4_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26043\,
            in1 => \N__36488\,
            in2 => \_gnd_net_\,
            in3 => \N__21477\,
            lcout => \dataRead7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38681\,
            ce => 'H',
            sr => \N__35707\
        );

    \QuadInstance0.Quad_9_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28565\,
            in1 => \N__33129\,
            in2 => \_gnd_net_\,
            in3 => \N__30117\,
            lcout => \dataRead0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38681\,
            ce => 'H',
            sr => \N__35707\
        );

    \QuadInstance1.un1_Quad_cry_0_c_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24196\,
            in2 => \N__30943\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \QuadInstance1.un1_Quad_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23890\,
            in2 => \N__23538\,
            in3 => \N__21636\,
            lcout => \QuadInstance1.Quad_RNO_0_0_1\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_0\,
            carryout => \QuadInstance1.un1_Quad_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30568\,
            in2 => \N__23676\,
            in3 => \N__21618\,
            lcout => \QuadInstance1.Quad_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_1\,
            carryout => \QuadInstance1.un1_Quad_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27874\,
            in2 => \N__23667\,
            in3 => \N__21603\,
            lcout => \QuadInstance1.Quad_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_2\,
            carryout => \QuadInstance1.un1_Quad_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23263\,
            in2 => \N__23241\,
            in3 => \N__21594\,
            lcout => \QuadInstance1.Quad_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_3\,
            carryout => \QuadInstance1.un1_Quad_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_5_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36817\,
            in2 => \N__23520\,
            in3 => \N__21582\,
            lcout => \QuadInstance1.Quad_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_4\,
            carryout => \QuadInstance1.un1_Quad_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_6_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25303\,
            in2 => \N__23529\,
            in3 => \N__21567\,
            lcout => \QuadInstance1.Quad_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_5\,
            carryout => \QuadInstance1.un1_Quad_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_7_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25567\,
            in2 => \N__23685\,
            in3 => \N__21555\,
            lcout => \QuadInstance1.Quad_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_6\,
            carryout => \QuadInstance1.un1_Quad_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_8_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37012\,
            in2 => \N__23634\,
            in3 => \N__21690\,
            lcout => \QuadInstance1.Quad_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \QuadInstance1.un1_Quad_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_9_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25531\,
            in2 => \N__23481\,
            in3 => \N__21687\,
            lcout => \QuadInstance1.Quad_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_8\,
            carryout => \QuadInstance1.un1_Quad_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_10_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35050\,
            in2 => \N__23472\,
            in3 => \N__21678\,
            lcout => \QuadInstance1.Quad_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_9\,
            carryout => \QuadInstance1.un1_Quad_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_11_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23362\,
            in2 => \N__23340\,
            in3 => \N__21666\,
            lcout => \QuadInstance1.Quad_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_10\,
            carryout => \QuadInstance1.un1_Quad_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_12_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24121\,
            in2 => \N__23658\,
            in3 => \N__21663\,
            lcout => \QuadInstance1.Quad_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_11\,
            carryout => \QuadInstance1.un1_Quad_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_13_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23917\,
            in2 => \N__23649\,
            in3 => \N__21660\,
            lcout => \QuadInstance1.Quad_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_12\,
            carryout => \QuadInstance1.un1_Quad_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_14_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23640\,
            in2 => \N__28189\,
            in3 => \N__21651\,
            lcout => \QuadInstance1.Quad_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \QuadInstance1.un1_Quad_cry_13\,
            carryout => \QuadInstance1.un1_Quad_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_15_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__23547\,
            in1 => \N__24050\,
            in2 => \N__31896\,
            in3 => \N__21648\,
            lcout => \dataRead1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38664\,
            ce => 'H',
            sr => \N__35722\
        );

    \QuadInstance0.Quad_1_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31218\,
            in1 => \N__29892\,
            in2 => \_gnd_net_\,
            in3 => \N__33126\,
            lcout => \dataRead0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38652\,
            ce => 'H',
            sr => \N__35733\
        );

    \QuadInstance6.Quad_9_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22790\,
            in1 => \N__28528\,
            in2 => \_gnd_net_\,
            in3 => \N__22221\,
            lcout => \dataRead6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38652\,
            ce => 'H',
            sr => \N__35733\
        );

    \QuadInstance2.Quad_1_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31219\,
            in1 => \N__22209\,
            in2 => \_gnd_net_\,
            in3 => \N__22189\,
            lcout => \dataRead2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38652\,
            ce => 'H',
            sr => \N__35733\
        );

    \QuadInstance3.Quad_1_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22029\,
            in1 => \N__31220\,
            in2 => \_gnd_net_\,
            in3 => \N__22013\,
            lcout => \dataRead3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38652\,
            ce => 'H',
            sr => \N__35733\
        );

    \QuadInstance3.Quad_4_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22012\,
            in1 => \_gnd_net_\,
            in2 => \N__36483\,
            in3 => \N__21855\,
            lcout => \dataRead3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38652\,
            ce => 'H',
            sr => \N__35733\
        );

    \QuadInstance1.Quad_9_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24102\,
            in1 => \N__28527\,
            in2 => \_gnd_net_\,
            in3 => \N__21813\,
            lcout => \dataRead1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38652\,
            ce => 'H',
            sr => \N__35733\
        );

    \QuadInstance6.Quad_0_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__22753\,
            in1 => \N__22550\,
            in2 => \N__31434\,
            in3 => \N__30799\,
            lcout => \dataRead6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38652\,
            ce => 'H',
            sr => \N__35733\
        );

    \QuadInstance7.Quad_0_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__30769\,
            in1 => \N__31407\,
            in2 => \N__26042\,
            in3 => \N__21807\,
            lcout => \dataRead7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38652\,
            ce => 'H',
            sr => \N__35733\
        );

    \QuadInstance6.delayedCh_B_2_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22467\,
            lcout => \QuadInstance6.delayedCh_BZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNIGENB1_10_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__34610\,
            in1 => \N__22721\,
            in2 => \N__22632\,
            in3 => \N__22548\,
            lcout => \QuadInstance6.Quad_RNIGENB1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.delayedCh_A_2_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22863\,
            lcout => \QuadInstance6.delayedCh_AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.Quad_RNIJHNB1_13_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__22838\,
            in1 => \N__22722\,
            in2 => \N__22633\,
            in3 => \N__22549\,
            lcout => \QuadInstance6.Quad_RNIJHNB1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.delayedCh_B_1_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27108\,
            lcout => \QuadInstance6.delayedCh_BZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_3_11_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__22450\,
            in1 => \N__34870\,
            in2 => \N__34772\,
            in3 => \N__22418\,
            lcout => \OutReg_0_4_i_m3_i_m3_ns_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_2_12_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__24129\,
            in1 => \N__38138\,
            in2 => \N__22389\,
            in3 => \N__27624\,
            lcout => \OutReg_esr_RNO_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_3_12_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__28126\,
            in1 => \N__22359\,
            in2 => \N__22331\,
            in3 => \N__28012\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_1_12_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__22293\,
            in1 => \N__22263\,
            in2 => \N__22233\,
            in3 => \N__37742\,
            lcout => OPEN,
            ltout => \OutReg_esr_RNO_1Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_0_12_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37559\,
            in2 => \N__22230\,
            in3 => \N__22227\,
            lcout => OPEN,
            ltout => \OutReg_esr_RNO_0Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_12_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__22941\,
            in1 => \N__38951\,
            in2 => \N__22932\,
            in3 => \N__37388\,
            lcout => \OutRegZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38633\,
            ce => \N__37242\,
            sr => \N__37130\
        );

    \data_received_esr_13_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22922\,
            lcout => \data_receivedZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38620\,
            ce => \N__26182\,
            sr => \N__26152\
        );

    \data_received_esr_10_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24474\,
            lcout => \data_receivedZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38620\,
            ce => \N__26182\,
            sr => \N__26152\
        );

    \data_received_esr_12_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22874\,
            lcout => \data_receivedZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38620\,
            ce => \N__26182\,
            sr => \N__26152\
        );

    \data_received_esr_14_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22910\,
            lcout => \data_receivedZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38620\,
            ce => \N__26182\,
            sr => \N__26152\
        );

    \data_received_esr_11_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22886\,
            lcout => \data_receivedZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38620\,
            ce => \N__26182\,
            sr => \N__26152\
        );

    \data_received_esr_23_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33283\,
            lcout => \data_receivedZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38620\,
            ce => \N__26182\,
            sr => \N__26152\
        );

    \pwmWrite_3_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33759\,
            in1 => \N__33557\,
            in2 => \N__33468\,
            in3 => \N__23391\,
            lcout => \pwmWriteZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_esr_RNIMIH31_19_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__22994\,
            in1 => \N__37985\,
            in2 => \N__22980\,
            in3 => \N__39064\,
            lcout => \data_received_esr_RNIMIH31Z0Z_19\,
            ltout => \data_received_esr_RNIMIH31Z0Z_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_fast_3_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33761\,
            in1 => \N__33459\,
            in2 => \N__22998\,
            in3 => \N__33559\,
            lcout => \pwmWrite_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_esr_RNIBPOR_23_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__22978\,
            in1 => \N__37986\,
            in2 => \_gnd_net_\,
            in3 => \N__39066\,
            lcout => \N_870_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_esr_RNIMIH31_0_19_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__22993\,
            in1 => \N__37984\,
            in2 => \N__22979\,
            in3 => \N__39065\,
            lcout => \data_received_esr_RNIMIH31_0Z0Z_19\,
            ltout => \data_received_esr_RNIMIH31_0Z0Z_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_fast_2_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33760\,
            in1 => \N__33458\,
            in2 => \N__22962\,
            in3 => \N__33558\,
            lcout => \pwmWrite_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_0_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31382\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38599\,
            ce => \N__26958\,
            sr => \N__35764\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_13_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28677\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38592\,
            ce => \N__24539\,
            sr => \N__35770\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_5_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36332\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38592\,
            ce => \N__24539\,
            sr => \N__35770\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_8_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28943\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38592\,
            ce => \N__24539\,
            sr => \N__35770\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_11_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35994\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38592\,
            ce => \N__24539\,
            sr => \N__35770\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_12_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28823\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38592\,
            ce => \N__24539\,
            sr => \N__35770\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__23195\,
            in1 => \N__23145\,
            in2 => \N__23139\,
            in3 => \N__23174\,
            lcout => \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_14_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34394\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38581\,
            ce => \N__24558\,
            sr => \N__35774\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_15_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31857\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38581\,
            ce => \N__24558\,
            sr => \N__35774\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23130\,
            in1 => \N__23109\,
            in2 => \N__23103\,
            in3 => \N__23067\,
            lcout => \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_10_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36158\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38581\,
            ce => \N__24558\,
            sr => \N__35774\
        );

    \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__23061\,
            in1 => \N__23055\,
            in2 => \N__23034\,
            in3 => \N__23010\,
            lcout => \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_12_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28854\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38571\,
            ce => \N__26953\,
            sr => \N__35782\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_13_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28711\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38571\,
            ce => \N__26953\,
            sr => \N__35782\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_8_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28976\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38571\,
            ce => \N__26953\,
            sr => \N__35782\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_9_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28557\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38571\,
            ce => \N__26953\,
            sr => \N__35782\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_3_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32043\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38571\,
            ce => \N__26953\,
            sr => \N__35782\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__23208\,
            in1 => \N__24652\,
            in2 => \N__24834\,
            in3 => \N__23214\,
            lcout => \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.periodCounter_RNI3G5D_2_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24910\,
            in2 => \_gnd_net_\,
            in3 => \N__24694\,
            lcout => OPEN,
            ltout => \PWMInstance4.un1_periodCounter12_1_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.periodCounter_RNIDRK61_4_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__24745\,
            in1 => \N__24797\,
            in2 => \N__23217\,
            in3 => \N__24653\,
            lcout => \PWMInstance4.un1_periodCounter12_1_0_a2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_4_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36502\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38563\,
            ce => \N__26952\,
            sr => \N__35786\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_5_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36362\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38563\,
            ce => \N__26952\,
            sr => \N__35786\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24796\,
            in1 => \N__23331\,
            in2 => \N__24776\,
            in3 => \N__23202\,
            lcout => \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_10_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36159\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38563\,
            ce => \N__26952\,
            sr => \N__35786\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_11_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36014\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38563\,
            ce => \N__26952\,
            sr => \N__35786\
        );

    \QuadInstance2.delayedCh_B_0_LC_14_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance2.delayedCh_BZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.delayedCh_B_0_LC_14_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23295\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance4.delayedCh_BZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.delayedCh_A_0_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23280\,
            lcout => \QuadInstance4.delayedCh_AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.delayedCh_B_1_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27072\,
            lcout => \QuadInstance1.delayedCh_BZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.delayedCh_B_2_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23231\,
            lcout => \QuadInstance1.delayedCh_BZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.delayedCh_A_1_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32118\,
            lcout => \QuadInstance1.delayedCh_AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNIRK0O_4_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \N__23264\,
            in1 => \N__23580\,
            in2 => \N__24084\,
            in3 => \N__24180\,
            lcout => \QuadInstance1.Quad_RNIRK0OZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.delayedCh_A_RNIGDO2_2_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23502\,
            in1 => \N__23492\,
            in2 => \N__23511\,
            in3 => \N__23232\,
            lcout => \QuadInstance1.count_enable\,
            ltout => \QuadInstance1.count_enable_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNIOH0O_1_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__23898\,
            in1 => \N__24004\,
            in2 => \N__23541\,
            in3 => \N__23579\,
            lcout => \QuadInstance1.Quad_RNIOH0OZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNITM0O_6_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001010"
        )
    port map (
            in0 => \N__24181\,
            in1 => \N__24052\,
            in2 => \N__23610\,
            in3 => \N__25311\,
            lcout => \QuadInstance1.Quad_RNITM0OZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNISL0O_5_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \N__36827\,
            in1 => \N__23581\,
            in2 => \N__24085\,
            in3 => \N__24182\,
            lcout => \QuadInstance1.Quad_RNISL0OZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.delayedCh_A_2_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23493\,
            lcout => \QuadInstance1.delayedCh_AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38690\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.delayedCh_B_RNIM2H8_2_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__23501\,
            in1 => \N__34495\,
            in2 => \_gnd_net_\,
            in3 => \N__23491\,
            lcout => \QuadInstance1.un1_count_enable_i_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNI0Q0O_9_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__25545\,
            in1 => \N__24008\,
            in2 => \N__24198\,
            in3 => \N__23595\,
            lcout => \QuadInstance1.Quad_RNI0Q0OZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNI8P5D_10_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__24009\,
            in1 => \N__35061\,
            in2 => \N__23613\,
            in3 => \N__24178\,
            lcout => \QuadInstance1.Quad_RNI8P5DZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quadWrite_1_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33858\,
            in1 => \N__33656\,
            in2 => \N__33448\,
            in3 => \N__23448\,
            lcout => \quadWriteZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNI9Q5D_11_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__24010\,
            in1 => \N__23370\,
            in2 => \N__23614\,
            in3 => \N__24179\,
            lcout => \QuadInstance1.Quad_RNI9Q5DZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_3_5_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__34731\,
            in1 => \N__23734\,
            in2 => \N__34889\,
            in3 => \N__23710\,
            lcout => \OutReg_0_4_i_m3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNIUN0O_7_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__24007\,
            in1 => \N__25568\,
            in2 => \N__23612\,
            in3 => \N__24174\,
            lcout => \QuadInstance1.Quad_RNIUN0OZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNIPI0O_2_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__30569\,
            in1 => \N__24005\,
            in2 => \N__24197\,
            in3 => \N__23588\,
            lcout => \QuadInstance1.Quad_RNIPI0OZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNIQJ0O_3_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__24006\,
            in1 => \N__27878\,
            in2 => \N__23611\,
            in3 => \N__24173\,
            lcout => \QuadInstance1.Quad_RNIQJ0OZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNIAR5D_12_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__24200\,
            in1 => \N__23618\,
            in2 => \N__24128\,
            in3 => \N__24022\,
            lcout => \QuadInstance1.Quad_RNIAR5DZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNIBS5D_13_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001100"
        )
    port map (
            in0 => \N__24023\,
            in1 => \N__24201\,
            in2 => \N__23625\,
            in3 => \N__23918\,
            lcout => \QuadInstance1.Quad_RNIBS5DZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNICT5D_14_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \N__28190\,
            in1 => \N__23622\,
            in2 => \N__24209\,
            in3 => \N__24024\,
            lcout => \QuadInstance1.Quad_RNICT5DZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNIVO0O_8_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__24021\,
            in1 => \N__37013\,
            in2 => \N__23624\,
            in3 => \N__24199\,
            lcout => \QuadInstance1.Quad_RNIVO0OZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_RNO_0_15_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010011010"
        )
    port map (
            in0 => \N__24227\,
            in1 => \N__23623\,
            in2 => \N__24210\,
            in3 => \N__24025\,
            lcout => \QuadInstance1.un1_Quad_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.Quad_0_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__24027\,
            in1 => \N__31411\,
            in2 => \N__30947\,
            in3 => \N__24208\,
            lcout => \dataRead1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38674\,
            ce => 'H',
            sr => \N__35734\
        );

    \QuadInstance1.Quad_12_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28833\,
            in1 => \N__24028\,
            in2 => \_gnd_net_\,
            in3 => \N__24135\,
            lcout => \dataRead1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38674\,
            ce => 'H',
            sr => \N__35734\
        );

    \QuadInstance1.Quad_13_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24026\,
            in1 => \N__28715\,
            in2 => \_gnd_net_\,
            in3 => \N__23928\,
            lcout => \dataRead1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38674\,
            ce => 'H',
            sr => \N__35734\
        );

    \OutReg_ess_RNO_2_1_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__23897\,
            in1 => \N__23751\,
            in2 => \N__23868\,
            in3 => \N__32926\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_0_1_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37502\,
            in2 => \N__23838\,
            in3 => \N__23757\,
            lcout => \OutReg_ess_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_3_1_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__23827\,
            in1 => \N__34732\,
            in2 => \N__34884\,
            in3 => \N__23800\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_1_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__25834\,
            in1 => \N__23787\,
            in2 => \N__23760\,
            in3 => \N__32811\,
            lcout => \OutReg_ess_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_4_1_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__32716\,
            in1 => \N__28102\,
            in2 => \N__27996\,
            in3 => \N__27220\,
            lcout => \OutReg_0_5_i_m3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_fast_esr_2_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37504\,
            lcout => \data_received_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38665\,
            ce => \N__26178\,
            sr => \N__26156\
        );

    \data_received_2_rep1_esr_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37503\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \data_received_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38665\,
            ce => \N__26178\,
            sr => \N__26156\
        );

    \OutReg_ess_RNO_3_3_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__34733\,
            in1 => \N__24410\,
            in2 => \N__24374\,
            in3 => \N__34862\,
            lcout => \OutReg_0_4_i_m3_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_15_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__38946\,
            in1 => \N__37374\,
            in2 => \N__26205\,
            in3 => \N__37821\,
            lcout => \OutRegZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38653\,
            ce => \N__37245\,
            sr => \N__37135\
        );

    \OutReg_ess_RNO_3_15_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__24336\,
            in1 => \N__24315\,
            in2 => \N__28016\,
            in3 => \N__28101\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_15_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__24291\,
            in1 => \N__24269\,
            in2 => \N__24249\,
            in3 => \N__37708\,
            lcout => \OutReg_ess_RNO_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_2_15_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001010101"
        )
    port map (
            in0 => \N__25197\,
            in1 => \N__24246\,
            in2 => \N__24228\,
            in3 => \N__38114\,
            lcout => \OutReg_ess_RNO_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_esr_5_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34979\,
            lcout => \data_receivedZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38643\,
            ce => \N__26183\,
            sr => \N__26153\
        );

    \data_received_esr_7_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24437\,
            lcout => \data_receivedZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38643\,
            ce => \N__26183\,
            sr => \N__26153\
        );

    \data_received_esr_9_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24485\,
            lcout => \data_receivedZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38643\,
            ce => \N__26183\,
            sr => \N__26153\
        );

    \data_received_esr_22_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33842\,
            lcout => \data_receivedZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38643\,
            ce => \N__26183\,
            sr => \N__26153\
        );

    \data_received_esr_6_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24449\,
            lcout => \data_receivedZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38643\,
            ce => \N__26183\,
            sr => \N__26153\
        );

    \data_received_esr_8_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24425\,
            lcout => \data_receivedZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38643\,
            ce => \N__26183\,
            sr => \N__26153\
        );

    \dataWrite_2_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37712\,
            lcout => \dataWriteZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__24462\,
            sr => \_gnd_net_\
        );

    \dataWrite_3_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30638\,
            lcout => \dataWriteZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__24462\,
            sr => \_gnd_net_\
        );

    \dataWrite_4_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34978\,
            lcout => \dataWriteZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__24462\,
            sr => \_gnd_net_\
        );

    \dataWrite_5_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24450\,
            lcout => \dataWriteZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__24462\,
            sr => \_gnd_net_\
        );

    \dataWrite_6_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24438\,
            lcout => \dataWriteZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__24462\,
            sr => \_gnd_net_\
        );

    \dataWrite_7_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24426\,
            lcout => \dataWriteZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__24462\,
            sr => \_gnd_net_\
        );

    \dataWrite_8_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24486\,
            lcout => \dataWriteZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__24462\,
            sr => \_gnd_net_\
        );

    \dataWrite_9_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24473\,
            lcout => \dataWriteZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__24462\,
            sr => \_gnd_net_\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_11_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35974\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38621\,
            ce => \N__29290\,
            sr => \N__35765\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_8_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28912\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38621\,
            ce => \N__29290\,
            sr => \N__35765\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_5_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36284\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38621\,
            ce => \N__29290\,
            sr => \N__35765\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_10_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36157\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38621\,
            ce => \N__29290\,
            sr => \N__35765\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_3_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31985\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38621\,
            ce => \N__29290\,
            sr => \N__35765\
        );

    \PWMInstance3.out_RNO_0_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__24621\,
            in1 => \N__24604\,
            in2 => \N__26709\,
            in3 => \N__24589\,
            lcout => \PWMInstance3.un1_periodCounter12_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.clkCount_0_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000101"
        )
    port map (
            in0 => \N__24590\,
            in1 => \_gnd_net_\,
            in2 => \N__24611\,
            in3 => \N__24635\,
            lcout => \PWMInstance3.clkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38612\,
            ce => 'H',
            sr => \N__35771\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_ctle_15_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__35830\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24634\,
            lcout => \PWMInstance3.pwmWrite_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.clkCount_1_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000001010"
        )
    port map (
            in0 => \N__24591\,
            in1 => \_gnd_net_\,
            in2 => \N__24612\,
            in3 => \N__24636\,
            lcout => \PWMInstance3.clkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38612\,
            ce => 'H',
            sr => \N__35771\
        );

    \PWMInstance3.clkCount_RNI21FG_0_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__24620\,
            in1 => \N__24603\,
            in2 => \_gnd_net_\,
            in3 => \N__24588\,
            lcout => \PWMInstance3.periodCounter12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.periodCounter_RNI8K3C_16_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26705\,
            in2 => \_gnd_net_\,
            in3 => \N__29497\,
            lcout => OPEN,
            ltout => \PWMInstance3.un1_periodCounter12_1_0_a2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.periodCounter_RNIB2M81_1_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__29038\,
            in1 => \N__29170\,
            in2 => \N__24576\,
            in3 => \N__26428\,
            lcout => OPEN,
            ltout => \PWMInstance3.un1_periodCounter12_1_0_a2_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.periodCounter_RNI0E0J3_0_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28389\,
            in1 => \N__29067\,
            in2 => \N__24573\,
            in3 => \N__26457\,
            lcout => \PWMInstance3.out_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance6.PWMPulseWidthCount_esr_9_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28523\,
            lcout => \PWMInstance6.PWMPulseWidthCountZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38600\,
            ce => \N__24552\,
            sr => \N__35775\
        );

    \PWMInstance4.periodCounter_RNIRPSE_3_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26550\,
            in1 => \N__24832\,
            in2 => \N__24780\,
            in3 => \N__24673\,
            lcout => \PWMInstance4.un1_periodCounter12_1_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__24498\,
            in1 => \N__24492\,
            in2 => \N__24675\,
            in3 => \N__24695\,
            lcout => \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_2_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38593\,
            ce => \N__26954\,
            sr => \N__35783\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__24717\,
            in1 => \N__24723\,
            in2 => \N__26841\,
            in3 => \N__24915\,
            lcout => \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_14_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34395\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38593\,
            ce => \N__26954\,
            sr => \N__35783\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_15_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31858\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38593\,
            ce => \N__26954\,
            sr => \N__35783\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24711\,
            in1 => \N__24705\,
            in2 => \N__26688\,
            in3 => \N__24750\,
            lcout => \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.periodCounter_0_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26664\,
            in2 => \N__26856\,
            in3 => \N__26855\,
            lcout => \PWMInstance4.periodCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_0\,
            clk => \N__38582\,
            ce => 'H',
            sr => \N__35297\
        );

    \PWMInstance4.periodCounter_1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26813\,
            in2 => \_gnd_net_\,
            in3 => \N__24699\,
            lcout => \PWMInstance4.periodCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_0\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_1\,
            clk => \N__38582\,
            ce => 'H',
            sr => \N__35297\
        );

    \PWMInstance4.periodCounter_2_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24696\,
            in2 => \_gnd_net_\,
            in3 => \N__24678\,
            lcout => \PWMInstance4.periodCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_1\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_2\,
            clk => \N__38582\,
            ce => 'H',
            sr => \N__35297\
        );

    \PWMInstance4.periodCounter_3_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24674\,
            in2 => \_gnd_net_\,
            in3 => \N__24657\,
            lcout => \PWMInstance4.periodCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_2\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_3\,
            clk => \N__38582\,
            ce => 'H',
            sr => \N__35297\
        );

    \PWMInstance4.periodCounter_4_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24654\,
            in2 => \_gnd_net_\,
            in3 => \N__24639\,
            lcout => \PWMInstance4.periodCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_3\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_4\,
            clk => \N__38582\,
            ce => 'H',
            sr => \N__35297\
        );

    \PWMInstance4.periodCounter_5_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24833\,
            in2 => \_gnd_net_\,
            in3 => \N__24813\,
            lcout => \PWMInstance4.periodCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_4\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_5\,
            clk => \N__38582\,
            ce => 'H',
            sr => \N__35297\
        );

    \PWMInstance4.periodCounter_6_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26619\,
            in2 => \_gnd_net_\,
            in3 => \N__24810\,
            lcout => \PWMInstance4.periodCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_5\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_6\,
            clk => \N__38582\,
            ce => 'H',
            sr => \N__35297\
        );

    \PWMInstance4.periodCounter_7_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26749\,
            in1 => \N__26994\,
            in2 => \_gnd_net_\,
            in3 => \N__24807\,
            lcout => \PWMInstance4.periodCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_6\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_7\,
            clk => \N__38582\,
            ce => 'H',
            sr => \N__35297\
        );

    \PWMInstance4.periodCounter_8_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26567\,
            in2 => \_gnd_net_\,
            in3 => \N__24804\,
            lcout => \PWMInstance4.periodCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_8\,
            clk => \N__38572\,
            ce => 'H',
            sr => \N__35295\
        );

    \PWMInstance4.periodCounter_9_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26548\,
            in2 => \_gnd_net_\,
            in3 => \N__24801\,
            lcout => \PWMInstance4.periodCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_8\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_9\,
            clk => \N__38572\,
            ce => 'H',
            sr => \N__35295\
        );

    \PWMInstance4.periodCounter_10_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24798\,
            in2 => \_gnd_net_\,
            in3 => \N__24783\,
            lcout => \PWMInstance4.periodCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_9\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_10\,
            clk => \N__38572\,
            ce => 'H',
            sr => \N__35295\
        );

    \PWMInstance4.periodCounter_11_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26747\,
            in1 => \N__24775\,
            in2 => \_gnd_net_\,
            in3 => \N__24753\,
            lcout => \PWMInstance4.periodCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_10\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_11\,
            clk => \N__38572\,
            ce => 'H',
            sr => \N__35295\
        );

    \PWMInstance4.periodCounter_12_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26746\,
            in1 => \N__24749\,
            in2 => \_gnd_net_\,
            in3 => \N__24729\,
            lcout => \PWMInstance4.periodCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_11\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_12\,
            clk => \N__38572\,
            ce => 'H',
            sr => \N__35295\
        );

    \PWMInstance4.periodCounter_13_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26748\,
            in1 => \N__26683\,
            in2 => \_gnd_net_\,
            in3 => \N__24726\,
            lcout => \PWMInstance4.periodCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_12\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_13\,
            clk => \N__38572\,
            ce => 'H',
            sr => \N__35295\
        );

    \PWMInstance4.periodCounter_14_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24914\,
            in2 => \_gnd_net_\,
            in3 => \N__24894\,
            lcout => \PWMInstance4.periodCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_13\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_14\,
            clk => \N__38572\,
            ce => 'H',
            sr => \N__35295\
        );

    \PWMInstance4.periodCounter_15_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26834\,
            in2 => \_gnd_net_\,
            in3 => \N__24891\,
            lcout => \PWMInstance4.periodCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_periodCounter_2_cry_14\,
            carryout => \PWMInstance4.un1_periodCounter_2_cry_15\,
            clk => \N__38572\,
            ce => 'H',
            sr => \N__35295\
        );

    \PWMInstance4.periodCounter_16_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26750\,
            in1 => \N__27009\,
            in2 => \_gnd_net_\,
            in3 => \N__24888\,
            lcout => \PWMInstance4.periodCounterZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38564\,
            ce => 'H',
            sr => \N__35293\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_LC_15_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26637\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_1_0_\,
            carryout => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_LC_15_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24885\,
            in2 => \N__32544\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_0\,
            carryout => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_LC_15_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24867\,
            in2 => \N__32538\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_1\,
            carryout => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_LC_15_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26604\,
            in2 => \N__32542\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_2\,
            carryout => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_LC_15_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26517\,
            in2 => \N__32540\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_3\,
            carryout => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_LC_15_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24852\,
            in2 => \N__32543\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_4\,
            carryout => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_LC_15_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25020\,
            in2 => \N__32539\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_5\,
            carryout => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_LC_15_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25002\,
            in2 => \N__32541\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_6\,
            carryout => \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.out_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__24962\,
            in1 => \N__27021\,
            in2 => \N__26757\,
            in3 => \N__24984\,
            lcout => \PWM4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38717\,
            ce => 'H',
            sr => \N__35701\
        );

    \QuadInstance4.un1_Quad_cry_0_c_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27432\,
            in2 => \N__30284\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_3_0_\,
            carryout => \QuadInstance4.un1_Quad_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_1_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27221\,
            in2 => \N__27195\,
            in3 => \N__24939\,
            lcout => \QuadInstance4.Quad_RNO_0_3_1\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_0\,
            carryout => \QuadInstance4.un1_Quad_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_2_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27178\,
            in2 => \N__27231\,
            in3 => \N__24936\,
            lcout => \QuadInstance4.Quad_RNO_0_4_2\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_1\,
            carryout => \QuadInstance4.un1_Quad_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_3_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28043\,
            in2 => \N__27159\,
            in3 => \N__24933\,
            lcout => \QuadInstance4.Quad_RNO_0_4_3\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_2\,
            carryout => \QuadInstance4.un1_Quad_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_4_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27528\,
            in2 => \N__27498\,
            in3 => \N__24918\,
            lcout => \QuadInstance4.Quad_RNO_0_4_4\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_3\,
            carryout => \QuadInstance4.un1_Quad_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_5_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27053\,
            in2 => \N__27036\,
            in3 => \N__25062\,
            lcout => \QuadInstance4.Quad_RNO_0_4_5\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_4\,
            carryout => \QuadInstance4.un1_Quad_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_6_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25087\,
            in2 => \N__25158\,
            in3 => \N__25059\,
            lcout => \QuadInstance4.Quad_RNO_0_4_6\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_5\,
            carryout => \QuadInstance4.un1_Quad_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_7_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27648\,
            in2 => \N__25239\,
            in3 => \N__25056\,
            lcout => \QuadInstance4.Quad_RNO_0_4_7\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_6\,
            carryout => \QuadInstance4.un1_Quad_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_8_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27264\,
            in2 => \N__27285\,
            in3 => \N__25053\,
            lcout => \QuadInstance4.Quad_RNO_0_4_8\,
            ltout => OPEN,
            carryin => \bfn_15_4_0_\,
            carryout => \QuadInstance4.un1_Quad_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_9_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25348\,
            in2 => \N__25251\,
            in3 => \N__25035\,
            lcout => \QuadInstance4.Quad_RNO_0_4_9\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_8\,
            carryout => \QuadInstance4.un1_Quad_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_10_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32867\,
            in2 => \N__25146\,
            in3 => \N__25032\,
            lcout => \QuadInstance4.Quad_RNO_0_4_10\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_9\,
            carryout => \QuadInstance4.un1_Quad_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_11_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25108\,
            in2 => \N__25137\,
            in3 => \N__25029\,
            lcout => \QuadInstance4.Quad_RNO_0_4_11\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_10\,
            carryout => \QuadInstance4.un1_Quad_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_12_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27027\,
            in2 => \N__27603\,
            in3 => \N__25026\,
            lcout => \QuadInstance4.Quad_RNO_0_4_12\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_11\,
            carryout => \QuadInstance4.un1_Quad_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_13_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27569\,
            in2 => \N__27150\,
            in3 => \N__25023\,
            lcout => \QuadInstance4.Quad_RNO_0_4_13\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_12\,
            carryout => \QuadInstance4.un1_Quad_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNO_0_14_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27141\,
            in2 => \N__29969\,
            in3 => \N__25188\,
            lcout => \QuadInstance4.Quad_RNO_0_4_14\,
            ltout => OPEN,
            carryin => \QuadInstance4.un1_Quad_cry_13\,
            carryout => \QuadInstance4.un1_Quad_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_15_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__25185\,
            in1 => \N__29628\,
            in2 => \N__31916\,
            in3 => \N__25170\,
            lcout => \dataRead4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38705\,
            ce => 'H',
            sr => \N__35716\
        );

    \QuadInstance0.Quad_6_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31107\,
            in1 => \N__33120\,
            in2 => \_gnd_net_\,
            in3 => \N__30243\,
            lcout => \dataRead0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38697\,
            ce => 'H',
            sr => \N__35723\
        );

    \QuadInstance4.Quad_6_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31108\,
            in1 => \N__29604\,
            in2 => \_gnd_net_\,
            in3 => \N__25167\,
            lcout => \dataRead4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38697\,
            ce => 'H',
            sr => \N__35723\
        );

    \QuadInstance4.Quad_RNIL00S1_6_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__29600\,
            in1 => \N__27423\,
            in2 => \N__25089\,
            in3 => \N__27342\,
            lcout => \QuadInstance4.Quad_RNIL00S1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNI06TL1_10_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010000"
        )
    port map (
            in0 => \N__27343\,
            in1 => \N__32871\,
            in2 => \N__27444\,
            in3 => \N__29601\,
            lcout => \QuadInstance4.Quad_RNI06TL1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNI17TL1_11_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__29602\,
            in1 => \N__27344\,
            in2 => \N__25115\,
            in3 => \N__27427\,
            lcout => \QuadInstance4.Quad_RNI17TL1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_11_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29603\,
            in1 => \N__36012\,
            in2 => \_gnd_net_\,
            in3 => \N__25128\,
            lcout => \dataRead4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38697\,
            ce => 'H',
            sr => \N__35723\
        );

    \OutReg_esr_RNO_4_6_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__33970\,
            in1 => \N__28127\,
            in2 => \N__25088\,
            in3 => \N__27976\,
            lcout => OPEN,
            ltout => \OutReg_0_5_i_m3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_2_6_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__25310\,
            in1 => \N__25280\,
            in2 => \N__25254\,
            in3 => \N__38094\,
            lcout => \OutReg_esr_RNO_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quadWrite_4_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33856\,
            in1 => \N__33658\,
            in2 => \N__33447\,
            in3 => \N__33234\,
            lcout => \quadWriteZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNIO30S1_9_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__29599\,
            in1 => \N__25349\,
            in2 => \N__27353\,
            in3 => \N__27439\,
            lcout => \QuadInstance4.Quad_RNIO30S1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_fast_4_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33855\,
            in1 => \N__33657\,
            in2 => \N__33446\,
            in3 => \N__33233\,
            lcout => \pwmWrite_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNIM10S1_7_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__27644\,
            in1 => \N__29598\,
            in2 => \N__27451\,
            in3 => \N__27338\,
            lcout => \QuadInstance4.Quad_RNIM10S1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_4_15_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__25214\,
            in1 => \N__32908\,
            in2 => \N__32818\,
            in3 => \N__30581\,
            lcout => \OutReg_0_5_i_m3_ns_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_15_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101001011010"
        )
    port map (
            in0 => \N__30582\,
            in1 => \N__33111\,
            in2 => \N__34086\,
            in3 => \N__33944\,
            lcout => \QuadInstance0.un1_Quad_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_0_rep2_esr_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35086\,
            lcout => \data_received_0_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38683\,
            ce => \N__26179\,
            sr => \N__26157\
        );

    \QuadInstance0.Quad_RNIOMBH1_9_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__30161\,
            in1 => \N__33110\,
            in2 => \N__34085\,
            in3 => \N__33943\,
            lcout => \QuadInstance0.Quad_RNIOMBH1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_0_rep1_esr_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35085\,
            lcout => \data_received_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38683\,
            ce => \N__26179\,
            sr => \N__26157\
        );

    \data_received_fast_esr_0_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35088\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \data_received_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38683\,
            ce => \N__26179\,
            sr => \N__26157\
        );

    \data_received_esr_0_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35087\,
            lcout => \data_receivedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38683\,
            ce => \N__26179\,
            sr => \N__26157\
        );

    \data_received_esr_1_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38100\,
            lcout => \data_receivedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38683\,
            ce => \N__26179\,
            sr => \N__26157\
        );

    \OutReg_ess_RNO_2_9_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__25544\,
            in1 => \N__38095\,
            in2 => \N__25518\,
            in3 => \N__25317\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_0_9_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37505\,
            in2 => \N__25485\,
            in3 => \N__25356\,
            lcout => \OutReg_ess_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_3_9_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__34742\,
            in1 => \N__25482\,
            in2 => \N__25452\,
            in3 => \N__34863\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_9_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__25414\,
            in1 => \N__25391\,
            in2 => \N__25359\,
            in3 => \N__37701\,
            lcout => \OutReg_ess_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_4_9_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__32810\,
            in1 => \N__30157\,
            in2 => \N__25350\,
            in3 => \N__32922\,
            lcout => \OutReg_0_5_i_m3_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_2_rep2_esr_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37507\,
            lcout => \data_received_2_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38675\,
            ce => \N__26180\,
            sr => \N__26155\
        );

    \data_received_esr_2_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37506\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \data_receivedZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38675\,
            ce => \N__26180\,
            sr => \N__26155\
        );

    \QuadInstance4.Quad_13_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28703\,
            in1 => \N__29642\,
            in2 => \_gnd_net_\,
            in3 => \N__26130\,
            lcout => \dataRead4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38666\,
            ce => 'H',
            sr => \N__35752\
        );

    \QuadInstance7.Quad_13_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28704\,
            in1 => \N__26040\,
            in2 => \_gnd_net_\,
            in3 => \N__26121\,
            lcout => \dataRead7_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38666\,
            ce => 'H',
            sr => \N__35752\
        );

    \QuadInstance4.Quad_3_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32020\,
            in1 => \N__29643\,
            in2 => \_gnd_net_\,
            in3 => \N__26079\,
            lcout => \dataRead4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38666\,
            ce => 'H',
            sr => \N__35752\
        );

    \QuadInstance7.Quad_3_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32022\,
            in1 => \N__26041\,
            in2 => \_gnd_net_\,
            in3 => \N__26070\,
            lcout => \dataRead7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38666\,
            ce => 'H',
            sr => \N__35752\
        );

    \QuadInstance7.Quad_1_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26039\,
            in1 => \N__31256\,
            in2 => \_gnd_net_\,
            in3 => \N__25857\,
            lcout => \dataRead7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38666\,
            ce => 'H',
            sr => \N__35752\
        );

    \QuadInstance5.Quad_3_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32021\,
            in1 => \N__25801\,
            in2 => \_gnd_net_\,
            in3 => \N__25641\,
            lcout => \dataRead5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38666\,
            ce => 'H',
            sr => \N__35752\
        );

    \GB_BUFFER_RST_c_i_g_THRU_LUT4_0_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35828\,
            lcout => \GB_BUFFER_RST_c_i_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_2_7_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__38139\,
            in1 => \N__25608\,
            in2 => \N__25575\,
            in3 => \N__27669\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_2Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_0_7_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__37537\,
            in1 => \_gnd_net_\,
            in2 => \N__26382\,
            in3 => \N__26235\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_7_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__28314\,
            in1 => \N__38879\,
            in2 => \N__26379\,
            in3 => \N__37378\,
            lcout => \OutRegZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38654\,
            ce => \N__37241\,
            sr => \N__37129\
        );

    \OutReg_ess_RNO_3_7_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__26376\,
            in1 => \N__34883\,
            in2 => \N__26340\,
            in3 => \N__34762\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_7_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__26304\,
            in1 => \N__26270\,
            in2 => \N__26238\,
            in3 => \N__37744\,
            lcout => \OutReg_ess_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_9_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__37379\,
            in1 => \N__37263\,
            in2 => \N__38910\,
            in3 => \N__26229\,
            lcout => \OutRegZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38654\,
            ce => \N__37241\,
            sr => \N__37129\
        );

    \OutReg_esr_14_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__38937\,
            in1 => \N__37380\,
            in2 => \N__26220\,
            in3 => \N__28146\,
            lcout => \OutRegZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38644\,
            ce => \N__37246\,
            sr => \N__37132\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__26190\,
            in1 => \N__26401\,
            in2 => \N__28437\,
            in3 => \N__26451\,
            lcout => \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.periodCounter_RNI1D3C_2_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29154\,
            in2 => \_gnd_net_\,
            in3 => \N__28348\,
            lcout => OPEN,
            ltout => \PWMInstance3.un1_periodCounter12_1_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.periodCounter_RNI83NV_4_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26493\,
            in1 => \N__29109\,
            in2 => \N__26460\,
            in3 => \N__26402\,
            lcout => \PWMInstance3.un1_periodCounter12_1_0_a2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_4_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36438\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38635\,
            ce => \N__29298\,
            sr => \N__35772\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__26445\,
            in1 => \N__26492\,
            in2 => \N__28416\,
            in3 => \N__26439\,
            lcout => \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.periodCounter_0_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29055\,
            in2 => \N__26433\,
            in3 => \N__26432\,
            lcout => \PWMInstance3.periodCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_0\,
            clk => \N__38622\,
            ce => 'H',
            sr => \N__35305\
        );

    \PWMInstance3.periodCounter_1_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29039\,
            in2 => \_gnd_net_\,
            in3 => \N__26412\,
            lcout => \PWMInstance3.periodCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_0\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_1\,
            clk => \N__38622\,
            ce => 'H',
            sr => \N__35305\
        );

    \PWMInstance3.periodCounter_2_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28350\,
            in2 => \_gnd_net_\,
            in3 => \N__26409\,
            lcout => \PWMInstance3.periodCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_1\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_2\,
            clk => \N__38622\,
            ce => 'H',
            sr => \N__35305\
        );

    \PWMInstance3.periodCounter_3_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28367\,
            in2 => \_gnd_net_\,
            in3 => \N__26406\,
            lcout => \PWMInstance3.periodCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_2\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_3\,
            clk => \N__38622\,
            ce => 'H',
            sr => \N__35305\
        );

    \PWMInstance3.periodCounter_4_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26403\,
            in2 => \_gnd_net_\,
            in3 => \N__26388\,
            lcout => \PWMInstance3.periodCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_3\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_4\,
            clk => \N__38622\,
            ce => 'H',
            sr => \N__35305\
        );

    \PWMInstance3.periodCounter_5_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28436\,
            in2 => \_gnd_net_\,
            in3 => \N__26385\,
            lcout => \PWMInstance3.periodCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_4\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_5\,
            clk => \N__38622\,
            ce => 'H',
            sr => \N__35305\
        );

    \PWMInstance3.periodCounter_6_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29481\,
            in2 => \_gnd_net_\,
            in3 => \N__26505\,
            lcout => \PWMInstance3.periodCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_5\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_6\,
            clk => \N__38622\,
            ce => 'H',
            sr => \N__35305\
        );

    \PWMInstance3.periodCounter_7_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29765\,
            in1 => \N__29501\,
            in2 => \_gnd_net_\,
            in3 => \N__26502\,
            lcout => \PWMInstance3.periodCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_6\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_7\,
            clk => \N__38622\,
            ce => 'H',
            sr => \N__35305\
        );

    \PWMInstance3.periodCounter_8_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29261\,
            in2 => \_gnd_net_\,
            in3 => \N__26499\,
            lcout => \PWMInstance3.periodCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_8\,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__35302\
        );

    \PWMInstance3.periodCounter_9_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29243\,
            in2 => \_gnd_net_\,
            in3 => \N__26496\,
            lcout => \PWMInstance3.periodCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_8\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_9\,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__35302\
        );

    \PWMInstance3.periodCounter_10_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26491\,
            in2 => \_gnd_net_\,
            in3 => \N__26475\,
            lcout => \PWMInstance3.periodCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_9\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_10\,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__35302\
        );

    \PWMInstance3.periodCounter_11_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29766\,
            in1 => \N__28411\,
            in2 => \_gnd_net_\,
            in3 => \N__26472\,
            lcout => \PWMInstance3.periodCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_10\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_11\,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__35302\
        );

    \PWMInstance3.periodCounter_12_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29764\,
            in1 => \N__29108\,
            in2 => \_gnd_net_\,
            in3 => \N__26469\,
            lcout => \PWMInstance3.periodCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_11\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_12\,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__35302\
        );

    \PWMInstance3.periodCounter_13_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29767\,
            in1 => \N__29087\,
            in2 => \_gnd_net_\,
            in3 => \N__26466\,
            lcout => \PWMInstance3.periodCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_12\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_13\,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__35302\
        );

    \PWMInstance3.periodCounter_14_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29153\,
            in2 => \_gnd_net_\,
            in3 => \N__26463\,
            lcout => \PWMInstance3.periodCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_13\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_14\,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__35302\
        );

    \PWMInstance3.periodCounter_15_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29174\,
            in2 => \_gnd_net_\,
            in3 => \N__26715\,
            lcout => \PWMInstance3.periodCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_periodCounter_2_cry_14\,
            carryout => \PWMInstance3.un1_periodCounter_2_cry_15\,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__35302\
        );

    \PWMInstance3.periodCounter_16_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29771\,
            in1 => \N__26704\,
            in2 => \_gnd_net_\,
            in3 => \N__26712\,
            lcout => \PWMInstance3.periodCounterZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38601\,
            ce => 'H',
            sr => \N__35300\
        );

    \PWMInstance4.periodCounter_RNIQOSE_0_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__26618\,
            in1 => \N__26684\,
            in2 => \N__26568\,
            in3 => \N__26663\,
            lcout => \PWMInstance4.un1_periodCounter12_1_0_a2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__26662\,
            in1 => \N__26625\,
            in2 => \N__26814\,
            in3 => \N__26649\,
            lcout => \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_1_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31281\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38594\,
            ce => \N__26934\,
            sr => \N__35789\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__26617\,
            in1 => \N__26592\,
            in2 => \N__26586\,
            in3 => \N__26993\,
            lcout => \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_6_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31118\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38594\,
            ce => \N__26934\,
            sr => \N__35789\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_7_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29418\,
            lcout => \PWMInstance4.PWMPulseWidthCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38594\,
            ce => \N__26934\,
            sr => \N__35789\
        );

    \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__26577\,
            in1 => \N__26563\,
            in2 => \N__26549\,
            in3 => \N__26526\,
            lcout => \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.out_RNO_0_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__26869\,
            in1 => \N__26904\,
            in2 => \N__26889\,
            in3 => \N__27008\,
            lcout => \PWMInstance4.un1_periodCounter12_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.clkCount_0_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__26975\,
            in1 => \N__26887\,
            in2 => \_gnd_net_\,
            in3 => \N__26870\,
            lcout => \PWMInstance4.clkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38583\,
            ce => 'H',
            sr => \N__35793\
        );

    \PWMInstance4.periodCounter_RNIAN5D_16_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27007\,
            in2 => \_gnd_net_\,
            in3 => \N__26992\,
            lcout => \PWMInstance4.un1_periodCounter12_1_0_a2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.clkCount_1_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110001000"
        )
    port map (
            in0 => \N__26976\,
            in1 => \N__26888\,
            in2 => \_gnd_net_\,
            in3 => \N__26871\,
            lcout => \PWMInstance4.clkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38583\,
            ce => 'H',
            sr => \N__35793\
        );

    \PWMInstance4.PWMPulseWidthCount_esr_ctle_15_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35832\,
            in2 => \_gnd_net_\,
            in3 => \N__26974\,
            lcout => \PWMInstance4.pwmWrite_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.clkCount_RNI5QJC_0_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__26903\,
            in1 => \N__26883\,
            in2 => \_gnd_net_\,
            in3 => \N__26868\,
            lcout => \PWMInstance4.periodCounter12\,
            ltout => \PWMInstance4.periodCounter12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.periodCounter_RNII1V61_1_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26833\,
            in1 => \N__26812\,
            in2 => \N__26793\,
            in3 => \N__26790\,
            lcout => OPEN,
            ltout => \PWMInstance4.un1_periodCounter12_1_0_a2_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance4.periodCounter_RNIKFDB3_0_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26784\,
            in1 => \N__26775\,
            in2 => \N__26769\,
            in3 => \N__26766\,
            lcout => \PWMInstance4.out_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance6.delayedCh_B_0_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27120\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance6.delayedCh_BZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM4_obufLegalizeSB_DFF_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM4_obufLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.delayedCh_B_0_LC_16_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27084\,
            lcout => \QuadInstance1.delayedCh_BZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_4_5_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__27052\,
            in1 => \N__28008\,
            in2 => \N__28139\,
            in3 => \N__34114\,
            lcout => \OutReg_0_5_i_m3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_5_LC_16_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29633\,
            in1 => \N__36347\,
            in2 => \_gnd_net_\,
            in3 => \N__27060\,
            lcout => \dataRead4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38718\,
            ce => 'H',
            sr => \N__35717\
        );

    \QuadInstance4.Quad_RNIKVVR1_5_LC_16_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__27054\,
            in1 => \N__29629\,
            in2 => \N__27445\,
            in3 => \N__27351\,
            lcout => \QuadInstance4.Quad_RNIKVVR1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNI28TL1_12_LC_16_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000100"
        )
    port map (
            in0 => \N__27352\,
            in1 => \N__27431\,
            in2 => \N__29652\,
            in3 => \N__27599\,
            lcout => \QuadInstance4.Quad_RNI28TL1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_4_2_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__32650\,
            in1 => \N__28132\,
            in2 => \N__27180\,
            in3 => \N__27989\,
            lcout => \OutReg_0_5_i_m3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_2_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31585\,
            in1 => \N__33130\,
            in2 => \_gnd_net_\,
            in3 => \N__29877\,
            lcout => \dataRead0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38711\,
            ce => 'H',
            sr => \N__35724\
        );

    \QuadInstance4.delayedCh_A_RNIS1AU_2_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27459\,
            in1 => \N__27474\,
            in2 => \N__29907\,
            in3 => \N__27134\,
            lcout => \QuadInstance4.count_enable\,
            ltout => \QuadInstance4.count_enable_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNIHSVR1_2_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__27179\,
            in1 => \N__29622\,
            in2 => \N__27234\,
            in3 => \N__27331\,
            lcout => \QuadInstance4.Quad_RNIHSVR1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNIGRVR1_1_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__27222\,
            in1 => \N__29621\,
            in2 => \N__27440\,
            in3 => \N__27330\,
            lcout => \QuadInstance4.Quad_RNIGRVR1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_2_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29624\,
            in1 => \N__31586\,
            in2 => \_gnd_net_\,
            in3 => \N__27186\,
            lcout => \dataRead4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38711\,
            ce => 'H',
            sr => \N__35724\
        );

    \QuadInstance4.Quad_RNIITVR1_3_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__28044\,
            in1 => \N__29623\,
            in2 => \N__27441\,
            in3 => \N__27332\,
            lcout => \QuadInstance4.Quad_RNIITVR1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.delayedCh_B_2_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29906\,
            lcout => \QuadInstance4.delayedCh_BZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNI39TL1_13_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__29589\,
            in1 => \N__27570\,
            in2 => \N__27443\,
            in3 => \N__27346\,
            lcout => \QuadInstance4.Quad_RNI39TL1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNI4ATL1_14_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__27347\,
            in1 => \N__29590\,
            in2 => \N__29965\,
            in3 => \N__27422\,
            lcout => \QuadInstance4.Quad_RNI4ATL1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.delayedCh_B_RNISS9M_2_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34496\,
            in2 => \N__27135\,
            in3 => \N__27472\,
            lcout => \QuadInstance4.un1_count_enable_i_a2_0_1\,
            ltout => \QuadInstance4.un1_count_enable_i_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNIJUVR1_4_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__27527\,
            in1 => \N__29587\,
            in2 => \N__27501\,
            in3 => \N__27415\,
            lcout => \QuadInstance4.Quad_RNIJUVR1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.delayedCh_A_1_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27486\,
            lcout => \QuadInstance4.delayedCh_AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.delayedCh_A_2_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27473\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance4.delayedCh_AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.Quad_RNIN20S1_8_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__29588\,
            in1 => \N__27263\,
            in2 => \N__27442\,
            in3 => \N__27345\,
            lcout => \QuadInstance4.Quad_RNIN20S1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_4_8_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__30193\,
            in1 => \N__32835\,
            in2 => \N__27259\,
            in3 => \N__32945\,
            lcout => \OutReg_0_5_i_m3_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_8_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33102\,
            in1 => \N__28990\,
            in2 => \_gnd_net_\,
            in3 => \N__30171\,
            lcout => \dataRead0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38698\,
            ce => 'H',
            sr => \N__35740\
        );

    \QuadInstance4.Quad_8_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28991\,
            in1 => \_gnd_net_\,
            in2 => \N__27276\,
            in3 => \N__29619\,
            lcout => \dataRead4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38698\,
            ce => 'H',
            sr => \N__35740\
        );

    \QuadInstance0.Quad_RNINLBH1_8_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__33101\,
            in1 => \N__30194\,
            in2 => \N__34081\,
            in3 => \N__33942\,
            lcout => \QuadInstance0.Quad_RNINLBH1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNIMKBH1_7_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__30227\,
            in1 => \N__33100\,
            in2 => \N__33950\,
            in3 => \N__34061\,
            lcout => \QuadInstance0.Quad_RNIMKBH1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_4_7_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__32946\,
            in1 => \N__27640\,
            in2 => \N__32841\,
            in3 => \N__30226\,
            lcout => \OutReg_0_5_i_m3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_7_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29426\,
            in1 => \N__33103\,
            in2 => \_gnd_net_\,
            in3 => \N__30204\,
            lcout => \dataRead0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38698\,
            ce => 'H',
            sr => \N__35740\
        );

    \QuadInstance4.Quad_7_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29618\,
            in1 => \N__29427\,
            in2 => \_gnd_net_\,
            in3 => \N__27657\,
            lcout => \dataRead4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38698\,
            ce => 'H',
            sr => \N__35740\
        );

    \OutReg_esr_RNO_4_12_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__32910\,
            in1 => \N__30049\,
            in2 => \N__27595\,
            in3 => \N__32801\,
            lcout => \OutReg_0_5_i_m3_ns_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_12_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33115\,
            in1 => \N__28861\,
            in2 => \_gnd_net_\,
            in3 => \N__30024\,
            lcout => \dataRead0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38692\,
            ce => 'H',
            sr => \N__35748\
        );

    \QuadInstance4.Quad_12_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28862\,
            in1 => \N__29620\,
            in2 => \_gnd_net_\,
            in3 => \N__27612\,
            lcout => \dataRead4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38692\,
            ce => 'H',
            sr => \N__35748\
        );

    \QuadInstance0.Quad_RNI2N8Q1_12_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__33113\,
            in1 => \N__30053\,
            in2 => \N__34087\,
            in3 => \N__33945\,
            lcout => \QuadInstance0.Quad_RNI2N8Q1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNI1M8Q1_11_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \N__30099\,
            in1 => \N__33112\,
            in2 => \N__33951\,
            in3 => \N__34077\,
            lcout => \QuadInstance0.Quad_RNI1M8Q1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNI3O8Q1_13_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010110000"
        )
    port map (
            in0 => \N__33114\,
            in1 => \N__33949\,
            in2 => \N__34088\,
            in3 => \N__30013\,
            lcout => \QuadInstance0.Quad_RNI3O8Q1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_4_13_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__32909\,
            in1 => \N__27565\,
            in2 => \N__30015\,
            in3 => \N__32800\,
            lcout => \OutReg_0_5_i_m3_ns_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_13_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33116\,
            in1 => \N__28727\,
            in2 => \_gnd_net_\,
            in3 => \N__29988\,
            lcout => \dataRead0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38692\,
            ce => 'H',
            sr => \N__35748\
        );

    \OutReg_ess_RNO_4_3_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__28128\,
            in1 => \N__34217\,
            in2 => \N__28042\,
            in3 => \N__27977\,
            lcout => OPEN,
            ltout => \OutReg_0_5_i_m3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_2_3_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__27913\,
            in1 => \N__27879\,
            in2 => \N__27846\,
            in3 => \N__38096\,
            lcout => \OutReg_ess_RNO_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_3_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__27843\,
            in1 => \N__37702\,
            in2 => \N__27816\,
            in3 => \N__27780\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_0_3_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37511\,
            in2 => \N__27771\,
            in3 => \N__27768\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_3_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__30474\,
            in1 => \N__38947\,
            in2 => \N__27762\,
            in3 => \N__37385\,
            lcout => \OutRegZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38684\,
            ce => \N__37250\,
            sr => \N__37136\
        );

    \OutReg_ess_4_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__37386\,
            in1 => \N__27759\,
            in2 => \N__38952\,
            in3 => \N__27753\,
            lcout => \OutRegZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38684\,
            ce => \N__37250\,
            sr => \N__37136\
        );

    \OutReg_esr_RNO_1_6_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__27741\,
            in1 => \N__37703\,
            in2 => \N__27708\,
            in3 => \N__28233\,
            lcout => OPEN,
            ltout => \OutReg_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_0_6_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37521\,
            in2 => \N__28332\,
            in3 => \N__28329\,
            lcout => OPEN,
            ltout => \OutReg_esr_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_6_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__38933\,
            in1 => \N__36666\,
            in2 => \N__28317\,
            in3 => \N__37351\,
            lcout => \OutRegZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38676\,
            ce => \N__37244\,
            sr => \N__37131\
        );

    \OutReg_esr_RNO_3_6_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__28304\,
            in1 => \N__34895\,
            in2 => \N__28269\,
            in3 => \N__34761\,
            lcout => \OutReg_0_4_i_m3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_esr_RNIA81U_3_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30634\,
            in1 => \N__37512\,
            in2 => \N__38137\,
            in3 => \N__37704\,
            lcout => \OutReg_0_sqmuxa_0_a2_3_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwmWrite_2_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33850\,
            in1 => \N__33660\,
            in2 => \N__33463\,
            in3 => \N__33214\,
            lcout => \pwmWriteZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_4_14_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__34251\,
            in1 => \N__32830\,
            in2 => \N__29970\,
            in3 => \N__32947\,
            lcout => OPEN,
            ltout => \OutReg_0_5_i_m3_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_2_14_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__28227\,
            in1 => \N__28191\,
            in2 => \N__28161\,
            in3 => \N__38113\,
            lcout => OPEN,
            ltout => \OutReg_esr_RNO_2Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_0_14_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__37513\,
            in1 => \_gnd_net_\,
            in2 => \N__28158\,
            in3 => \N__28155\,
            lcout => \OutReg_esr_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_12_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28819\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38655\,
            ce => \N__35854\,
            sr => \N__35773\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_13_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28699\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38655\,
            ce => \N__35854\,
            sr => \N__35773\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_8_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28972\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38655\,
            ce => \N__35854\,
            sr => \N__35773\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_9_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28506\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38655\,
            ce => \N__35854\,
            sr => \N__35773\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_7_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29392\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38655\,
            ce => \N__35854\,
            sr => \N__35773\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_12_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28871\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38645\,
            ce => \N__29319\,
            sr => \N__35776\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_13_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28724\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38645\,
            ce => \N__29319\,
            sr => \N__35776\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_9_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28541\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38645\,
            ce => \N__29319\,
            sr => \N__35776\
        );

    \PWMInstance3.periodCounter_RNINK9L_3_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__29242\,
            in1 => \N__28435\,
            in2 => \N__28415\,
            in3 => \N__28366\,
            lcout => \PWMInstance3.un1_periodCounter12_1_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__28380\,
            in1 => \N__29181\,
            in2 => \N__28368\,
            in3 => \N__28349\,
            lcout => \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_2_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31583\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38636\,
            ce => \N__29308\,
            sr => \N__35784\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__29133\,
            in1 => \N__29127\,
            in2 => \N__29175\,
            in3 => \N__29152\,
            lcout => \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_14_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34401\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38636\,
            ce => \N__29308\,
            sr => \N__35784\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_15_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31903\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38636\,
            ce => \N__29308\,
            sr => \N__35784\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__29121\,
            in1 => \N__29115\,
            in2 => \N__29088\,
            in3 => \N__29107\,
            lcout => \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.periodCounter_RNIMJ9L_0_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__29054\,
            in1 => \N__29083\,
            in2 => \N__29262\,
            in3 => \N__29479\,
            lcout => \PWMInstance3.un1_periodCounter12_1_0_a2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__29013\,
            in1 => \N__29053\,
            in2 => \N__29040\,
            in3 => \N__29019\,
            lcout => \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_0_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31412\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38623\,
            ce => \N__29318\,
            sr => \N__35787\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_1_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31280\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38623\,
            ce => \N__29318\,
            sr => \N__35787\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__29325\,
            in1 => \N__29466\,
            in2 => \N__29502\,
            in3 => \N__29480\,
            lcout => \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_6_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31094\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38623\,
            ce => \N__29318\,
            sr => \N__35787\
        );

    \PWMInstance3.PWMPulseWidthCount_esr_7_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance3.PWMPulseWidthCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38623\,
            ce => \N__29318\,
            sr => \N__35787\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__29274\,
            in1 => \N__29257\,
            in2 => \N__29244\,
            in3 => \N__29223\,
            lcout => \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29214\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29208\,
            in2 => \N__32579\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_0\,
            carryout => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29199\,
            in2 => \N__32573\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_1\,
            carryout => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29187\,
            in2 => \N__32577\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_2\,
            carryout => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29820\,
            in2 => \N__32575\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_3\,
            carryout => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29814\,
            in2 => \N__32578\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_4\,
            carryout => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29805\,
            in2 => \N__32574\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_5\,
            carryout => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29796\,
            in2 => \N__32576\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_6\,
            carryout => \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance3.out_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__29717\,
            in1 => \N__29787\,
            in2 => \N__29775\,
            in3 => \N__29730\,
            lcout => \PWM3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38602\,
            ce => 'H',
            sr => \N__35794\
        );

    \QuadInstance7.delayedCh_A_0_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29706\,
            lcout => \QuadInstance7.delayedCh_AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_5_LC_17_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36346\,
            in1 => \N__33109\,
            in2 => \_gnd_net_\,
            in3 => \N__29832\,
            lcout => \dataRead0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38722\,
            ce => 'H',
            sr => \N__35725\
        );

    \QuadInstance4.Quad_10_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__36165\,
            in1 => \_gnd_net_\,
            in2 => \N__29676\,
            in3 => \N__29661\,
            lcout => \dataRead4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38719\,
            ce => 'H',
            sr => \N__35735\
        );

    \QuadInstance4.Quad_14_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34416\,
            in1 => \N__29660\,
            in2 => \_gnd_net_\,
            in3 => \N__29979\,
            lcout => \dataRead4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38719\,
            ce => 'H',
            sr => \N__35735\
        );

    \QuadInstance0.delayedCh_B_1_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29934\,
            lcout => \QuadInstance0.delayedCh_BZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance4.delayedCh_B_1_LC_17_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29919\,
            lcout => \QuadInstance4.delayedCh_BZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.un1_Quad_cry_0_c_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34046\,
            in2 => \N__30317\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_6_0_\,
            carryout => \QuadInstance0.un1_Quad_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_1_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32729\,
            in2 => \N__32697\,
            in3 => \N__29880\,
            lcout => \QuadInstance0.Quad_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_0\,
            carryout => \QuadInstance0.un1_Quad_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_2_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32657\,
            in2 => \N__32637\,
            in3 => \N__29868\,
            lcout => \QuadInstance0.Quad_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_1\,
            carryout => \QuadInstance0.un1_Quad_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_3_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34176\,
            in2 => \N__34218\,
            in3 => \N__29850\,
            lcout => \QuadInstance0.Quad_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_2\,
            carryout => \QuadInstance0.un1_Quad_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_4_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34163\,
            in2 => \N__34134\,
            in3 => \N__29835\,
            lcout => \QuadInstance0.Quad_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_3\,
            carryout => \QuadInstance0.un1_Quad_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_5_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34121\,
            in2 => \N__34098\,
            in3 => \N__29823\,
            lcout => \QuadInstance0.Quad_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_4\,
            carryout => \QuadInstance0.un1_Quad_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_6_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33980\,
            in2 => \N__33867\,
            in3 => \N__30231\,
            lcout => \QuadInstance0.Quad_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_5\,
            carryout => \QuadInstance0.un1_Quad_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_7_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30228\,
            in2 => \N__30213\,
            in3 => \N__30198\,
            lcout => \QuadInstance0.Quad_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_6\,
            carryout => \QuadInstance0.un1_Quad_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_8_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30195\,
            in2 => \N__30180\,
            in3 => \N__30165\,
            lcout => \QuadInstance0.Quad_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => \QuadInstance0.un1_Quad_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_9_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30162\,
            in2 => \N__30129\,
            in3 => \N__30105\,
            lcout => \QuadInstance0.Quad_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_8\,
            carryout => \QuadInstance0.un1_Quad_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_10_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32687\,
            in2 => \N__32670\,
            in3 => \N__30102\,
            lcout => \QuadInstance0.Quad_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_9\,
            carryout => \QuadInstance0.un1_Quad_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_11_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30098\,
            in2 => \N__30075\,
            in3 => \N__30057\,
            lcout => \QuadInstance0.Quad_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_10\,
            carryout => \QuadInstance0.un1_Quad_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_12_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30054\,
            in2 => \N__30033\,
            in3 => \N__30018\,
            lcout => \QuadInstance0.Quad_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_11\,
            carryout => \QuadInstance0.un1_Quad_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_13_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30014\,
            in2 => \N__29997\,
            in3 => \N__29982\,
            lcout => \QuadInstance0.Quad_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_12\,
            carryout => \QuadInstance0.un1_Quad_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNO_0_14_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34224\,
            in2 => \N__34250\,
            in3 => \N__30597\,
            lcout => \QuadInstance0.Quad_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \QuadInstance0.un1_Quad_cry_13\,
            carryout => \QuadInstance0.un1_Quad_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_15_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__30594\,
            in1 => \N__33044\,
            in2 => \N__31917\,
            in3 => \N__30585\,
            lcout => \dataRead0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38699\,
            ce => 'H',
            sr => \N__35753\
        );

    \OutReg_esr_RNO_2_2_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__30570\,
            in1 => \N__38154\,
            in2 => \N__30534\,
            in3 => \N__30492\,
            lcout => OPEN,
            ltout => \OutReg_esr_RNO_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_0_2_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37557\,
            in2 => \N__30480\,
            in3 => \N__30324\,
            lcout => OPEN,
            ltout => \OutReg_esr_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_2_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__37332\,
            in1 => \N__30717\,
            in2 => \N__30477\,
            in3 => \N__38932\,
            lcout => \OutRegZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38693\,
            ce => \N__37224\,
            sr => \N__37115\
        );

    \OutReg_esr_RNO_3_2_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__30460\,
            in1 => \N__34885\,
            in2 => \N__30426\,
            in3 => \N__34764\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_1_2_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__30387\,
            in1 => \N__30353\,
            in2 => \N__30327\,
            in3 => \N__32831\,
            lcout => \OutReg_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_4_0_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__37763\,
            in1 => \N__30318\,
            in2 => \N__30285\,
            in3 => \N__38155\,
            lcout => OPEN,
            ltout => \OutReg_0_5_i_m3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_0_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__38156\,
            in1 => \N__30951\,
            in2 => \N__30918\,
            in3 => \N__30915\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_0_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__30747\,
            in1 => \N__34944\,
            in2 => \N__30885\,
            in3 => \N__37562\,
            lcout => \OutRegZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38685\,
            ce => \N__37210\,
            sr => \N__37128\
        );

    \OutReg_ess_RNO_3_0_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__30882\,
            in1 => \N__37761\,
            in2 => \N__30849\,
            in3 => \N__32949\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_0_0_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__37762\,
            in1 => \N__30809\,
            in2 => \N__30780\,
            in3 => \N__30777\,
            lcout => \OutReg_ess_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_1_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__37323\,
            in1 => \N__38913\,
            in2 => \N__30741\,
            in3 => \N__30729\,
            lcout => \OutRegZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38685\,
            ce => \N__37210\,
            sr => \N__37128\
        );

    \OutReg_esr_RNO_3_8_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__30710\,
            in1 => \N__34894\,
            in2 => \N__30675\,
            in3 => \N__34771\,
            lcout => \OutReg_0_4_i_m3_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_esr_RNI7L871_3_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__37313\,
            in1 => \N__38878\,
            in2 => \N__30642\,
            in3 => \N__39078\,
            lcout => OPEN,
            ltout => \data_received_esr_RNI7L871Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_esr_RNIKE1M2_3_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30600\,
            in3 => \N__37060\,
            lcout => \N_863_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_received_esr_RNIDPOE1_3_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__38877\,
            in1 => \N__37312\,
            in2 => \_gnd_net_\,
            in3 => \N__31446\,
            lcout => \OutReg_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.periodCounter_RNIIEMR_13_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34550\,
            in1 => \N__35422\,
            in2 => \N__35154\,
            in3 => \N__35107\,
            lcout => \PWMInstance2.un1_periodCounter12_1_0_a2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__31137\,
            in1 => \N__34549\,
            in2 => \N__35208\,
            in3 => \N__31287\,
            lcout => \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_0_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31437\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38668\,
            ce => \N__35861\,
            sr => \N__35777\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_1_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31240\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38668\,
            ce => \N__35861\,
            sr => \N__35777\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__31131\,
            in1 => \N__30969\,
            in2 => \N__35153\,
            in3 => \N__35129\,
            lcout => \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_6_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31063\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38668\,
            ce => \N__35861\,
            sr => \N__35777\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__30963\,
            in1 => \N__35455\,
            in2 => \N__35109\,
            in3 => \N__30957\,
            lcout => \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.out_RNO_0_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__31677\,
            in1 => \N__31657\,
            in2 => \N__35334\,
            in3 => \N__31642\,
            lcout => \PWMInstance2.un1_periodCounter12_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.clkCount_0_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000101"
        )
    port map (
            in0 => \N__31643\,
            in1 => \_gnd_net_\,
            in2 => \N__31664\,
            in3 => \N__31691\,
            lcout => \PWMInstance2.clkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38656\,
            ce => 'H',
            sr => \N__35785\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_ctle_15_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__31690\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35831\,
            lcout => \PWMInstance2.pwmWrite_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.clkCount_1_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000001010"
        )
    port map (
            in0 => \N__31644\,
            in1 => \_gnd_net_\,
            in2 => \N__31665\,
            in3 => \N__31692\,
            lcout => \PWMInstance2.clkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38656\,
            ce => 'H',
            sr => \N__35785\
        );

    \PWMInstance2.clkCount_RNIV7AK_0_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__31676\,
            in1 => \N__31656\,
            in2 => \_gnd_net_\,
            in3 => \N__31641\,
            lcout => \PWMInstance2.periodCounter12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.periodCounter_RNI6H1B_16_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35329\,
            in2 => \_gnd_net_\,
            in3 => \N__35128\,
            lcout => OPEN,
            ltout => \PWMInstance2.un1_periodCounter12_1_0_a2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.periodCounter_RNI43DA1_15_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__35395\,
            in1 => \N__35206\,
            in2 => \N__31629\,
            in3 => \N__34567\,
            lcout => OPEN,
            ltout => \PWMInstance2.un1_periodCounter12_1_0_a2_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.periodCounter_RNICCJQ3_10_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36534\,
            in1 => \N__31626\,
            in2 => \N__31620\,
            in3 => \N__31617\,
            lcout => \PWMInstance2.out_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.periodCounter_RNIJFMR_11_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__35180\,
            in1 => \N__35456\,
            in2 => \N__36200\,
            in3 => \N__35237\,
            lcout => \PWMInstance2.un1_periodCounter12_1_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__31935\,
            in1 => \N__35181\,
            in2 => \N__31455\,
            in3 => \N__36597\,
            lcout => \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_2_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31584\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38646\,
            ce => \N__35853\,
            sr => \N__35788\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_3_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32033\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38646\,
            ce => \N__35853\,
            sr => \N__35788\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__31737\,
            in1 => \N__31929\,
            in2 => \N__35400\,
            in3 => \N__36616\,
            lcout => \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_14_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34400\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38646\,
            ce => \N__35853\,
            sr => \N__35788\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_15_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31904\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38646\,
            ce => \N__35853\,
            sr => \N__35788\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__31731\,
            in1 => \N__31719\,
            in2 => \N__35427\,
            in3 => \N__36556\,
            lcout => \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31710\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32390\,
            in2 => \N__31701\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_0\,
            carryout => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35214\,
            in2 => \N__32494\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_1\,
            carryout => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32383\,
            in2 => \N__32619\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_2\,
            carryout => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32607\,
            in2 => \N__32496\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_3\,
            carryout => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36174\,
            in2 => \N__32518\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_4\,
            carryout => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32598\,
            in2 => \N__32495\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_5\,
            carryout => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32382\,
            in2 => \N__32172\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_6\,
            carryout => \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.out_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__32141\,
            in1 => \N__32163\,
            in2 => \N__35376\,
            in3 => \N__32154\,
            lcout => \PWM2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38624\,
            ce => 'H',
            sr => \N__35795\
        );

    \MOSIr_0_LC_18_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32130\,
            lcout => \MOSIrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38723\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance1.delayedCh_A_0_LC_18_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32124\,
            lcout => \QuadInstance1.delayedCh_AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38723\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.delayedCh_A_1_LC_18_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32106\,
            lcout => \QuadInstance0.delayedCh_AZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.delayedCh_A_2_LC_18_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34534\,
            lcout => \QuadInstance0.delayedCh_AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.delayedCh_B_2_LC_18_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32751\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \QuadInstance0.delayedCh_BZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_4_10_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__32944\,
            in1 => \N__32866\,
            in2 => \N__32840\,
            in3 => \N__32683\,
            lcout => \OutReg_0_5_i_m3_ns_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_10_LC_18_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33048\,
            in1 => \_gnd_net_\,
            in2 => \N__36164\,
            in3 => \N__32757\,
            lcout => \dataRead0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38713\,
            ce => 'H',
            sr => \N__35754\
        );

    \QuadInstance0.delayedCh_A_RNICHIP_2_LC_18_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32627\,
            in1 => \N__32750\,
            in2 => \N__34536\,
            in3 => \N__32739\,
            lcout => \QuadInstance0.count_enable\,
            ltout => \QuadInstance0.count_enable_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNIGEBH1_1_LC_18_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__32733\,
            in1 => \N__33045\,
            in2 => \N__32700\,
            in3 => \N__33903\,
            lcout => \QuadInstance0.Quad_RNIGEBH1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNI0L8Q1_10_LC_18_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__33047\,
            in1 => \N__33924\,
            in2 => \N__32688\,
            in3 => \N__34028\,
            lcout => \QuadInstance0.Quad_RNI0L8Q1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNIHFBH1_2_LC_18_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__32661\,
            in1 => \N__33046\,
            in2 => \N__34048\,
            in3 => \N__33904\,
            lcout => \QuadInstance0.Quad_RNIHFBH1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.delayedCh_B_RNIK4UJ_2_LC_18_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__32628\,
            in1 => \_gnd_net_\,
            in2 => \N__34535\,
            in3 => \N__34511\,
            lcout => \QuadInstance0.un1_count_enable_i_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_14_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34415\,
            in1 => \_gnd_net_\,
            in2 => \N__33053\,
            in3 => \N__34257\,
            lcout => \dataRead0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38707\,
            ce => 'H',
            sr => \N__35758\
        );

    \QuadInstance0.Quad_RNI4P8Q1_14_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100010"
        )
    port map (
            in0 => \N__34047\,
            in1 => \N__33913\,
            in2 => \N__33052\,
            in3 => \N__34249\,
            lcout => \QuadInstance0.Quad_RNI4P8Q1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNIIGBH1_3_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001010"
        )
    port map (
            in0 => \N__34030\,
            in1 => \N__34207\,
            in2 => \N__33925\,
            in3 => \N__33012\,
            lcout => \QuadInstance0.Quad_RNIIGBH1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNIJHBH1_4_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__33014\,
            in1 => \N__34029\,
            in2 => \N__34170\,
            in3 => \N__33905\,
            lcout => \QuadInstance0.Quad_RNIJHBH1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNIKIBH1_5_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001010"
        )
    port map (
            in0 => \N__34032\,
            in1 => \N__34125\,
            in2 => \N__33926\,
            in3 => \N__33013\,
            lcout => \QuadInstance0.Quad_RNIKIBH1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \QuadInstance0.Quad_RNILJBH1_6_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__33015\,
            in1 => \N__34031\,
            in2 => \N__33984\,
            in3 => \N__33909\,
            lcout => \QuadInstance0.Quad_RNILJBH1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quadWrite_0_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33851\,
            in1 => \N__33619\,
            in2 => \N__33400\,
            in3 => \N__33232\,
            lcout => \quadWriteZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \MOSIr_1_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32958\,
            lcout => \MOSIrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_2_10_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__35060\,
            in1 => \N__38159\,
            in2 => \N__35025\,
            in3 => \N__34989\,
            lcout => \OutReg_esr_RNO_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_RNI5AMB_0_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__37961\,
            in1 => \N__37886\,
            in2 => \N__34980\,
            in3 => \N__37812\,
            lcout => \un1_OutReg51_4_0_i_o3_2\,
            ltout => \un1_OutReg51_4_0_i_o3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_2_0_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34947\,
            in3 => \N__38912\,
            lcout => \OutReg_21_m_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_0_10_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37561\,
            in1 => \N__34578\,
            in2 => \_gnd_net_\,
            in3 => \N__34938\,
            lcout => \OutReg_esr_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_10_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__38900\,
            in1 => \N__37322\,
            in2 => \N__34932\,
            in3 => \N__34917\,
            lcout => \OutRegZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38686\,
            ce => \N__37211\,
            sr => \N__37099\
        );

    \OutReg_esr_RNO_3_10_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__34893\,
            in1 => \N__34802\,
            in2 => \N__34773\,
            in3 => \N__34683\,
            lcout => OPEN,
            ltout => \OutReg_0_4_i_m3_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_1_10_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__34649\,
            in1 => \N__34614\,
            in2 => \N__34581\,
            in3 => \N__37743\,
            lcout => \OutReg_esr_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.periodCounter_0_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34551\,
            in2 => \N__34572\,
            in3 => \N__34571\,
            lcout => \PWMInstance2.periodCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_0\,
            clk => \N__38677\,
            ce => 'H',
            sr => \N__35310\
        );

    \PWMInstance2.periodCounter_1_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35207\,
            in2 => \_gnd_net_\,
            in3 => \N__35187\,
            lcout => \PWMInstance2.periodCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_0\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_1\,
            clk => \N__38677\,
            ce => 'H',
            sr => \N__35310\
        );

    \PWMInstance2.periodCounter_2_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36595\,
            in2 => \_gnd_net_\,
            in3 => \N__35184\,
            lcout => \PWMInstance2.periodCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_1\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_2\,
            clk => \N__38677\,
            ce => 'H',
            sr => \N__35310\
        );

    \PWMInstance2.periodCounter_3_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35179\,
            in2 => \_gnd_net_\,
            in3 => \N__35163\,
            lcout => \PWMInstance2.periodCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_2\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_3\,
            clk => \N__38677\,
            ce => 'H',
            sr => \N__35310\
        );

    \PWMInstance2.periodCounter_4_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36574\,
            in2 => \_gnd_net_\,
            in3 => \N__35160\,
            lcout => \PWMInstance2.periodCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_3\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_4\,
            clk => \N__38677\,
            ce => 'H',
            sr => \N__35310\
        );

    \PWMInstance2.periodCounter_5_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35233\,
            in2 => \_gnd_net_\,
            in3 => \N__35157\,
            lcout => \PWMInstance2.periodCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_4\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_5\,
            clk => \N__38677\,
            ce => 'H',
            sr => \N__35310\
        );

    \PWMInstance2.periodCounter_6_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35152\,
            in2 => \_gnd_net_\,
            in3 => \N__35133\,
            lcout => \PWMInstance2.periodCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_5\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_6\,
            clk => \N__38677\,
            ce => 'H',
            sr => \N__35310\
        );

    \PWMInstance2.periodCounter_7_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35371\,
            in1 => \N__35130\,
            in2 => \_gnd_net_\,
            in3 => \N__35112\,
            lcout => \PWMInstance2.periodCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_6\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_7\,
            clk => \N__38677\,
            ce => 'H',
            sr => \N__35310\
        );

    \PWMInstance2.periodCounter_8_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35108\,
            in2 => \_gnd_net_\,
            in3 => \N__35091\,
            lcout => \PWMInstance2.periodCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_8\,
            clk => \N__38669\,
            ce => 'H',
            sr => \N__35309\
        );

    \PWMInstance2.periodCounter_9_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35457\,
            in2 => \_gnd_net_\,
            in3 => \N__35439\,
            lcout => \PWMInstance2.periodCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_8\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_9\,
            clk => \N__38669\,
            ce => 'H',
            sr => \N__35309\
        );

    \PWMInstance2.periodCounter_10_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36217\,
            in2 => \_gnd_net_\,
            in3 => \N__35436\,
            lcout => \PWMInstance2.periodCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_9\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_10\,
            clk => \N__38669\,
            ce => 'H',
            sr => \N__35309\
        );

    \PWMInstance2.periodCounter_11_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35369\,
            in1 => \N__36196\,
            in2 => \_gnd_net_\,
            in3 => \N__35433\,
            lcout => \PWMInstance2.periodCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_10\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_11\,
            clk => \N__38669\,
            ce => 'H',
            sr => \N__35309\
        );

    \PWMInstance2.periodCounter_12_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35368\,
            in1 => \N__36557\,
            in2 => \_gnd_net_\,
            in3 => \N__35430\,
            lcout => \PWMInstance2.periodCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_11\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_12\,
            clk => \N__38669\,
            ce => 'H',
            sr => \N__35309\
        );

    \PWMInstance2.periodCounter_13_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35370\,
            in1 => \N__35426\,
            in2 => \_gnd_net_\,
            in3 => \N__35406\,
            lcout => \PWMInstance2.periodCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_12\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_13\,
            clk => \N__38669\,
            ce => 'H',
            sr => \N__35309\
        );

    \PWMInstance2.periodCounter_14_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36617\,
            in2 => \_gnd_net_\,
            in3 => \N__35403\,
            lcout => \PWMInstance2.periodCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_13\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_14\,
            clk => \N__38669\,
            ce => 'H',
            sr => \N__35309\
        );

    \PWMInstance2.periodCounter_15_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35399\,
            in2 => \_gnd_net_\,
            in3 => \N__35379\,
            lcout => \PWMInstance2.periodCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \PWMInstance2.un1_periodCounter_2_cry_14\,
            carryout => \PWMInstance2.un1_periodCounter_2_cry_15\,
            clk => \N__38669\,
            ce => 'H',
            sr => \N__35309\
        );

    \PWMInstance2.periodCounter_16_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35372\,
            in1 => \N__35333\,
            in2 => \_gnd_net_\,
            in3 => \N__35337\,
            lcout => \PWMInstance2.periodCounterZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38657\,
            ce => 'H',
            sr => \N__35308\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36575\,
            in1 => \N__36225\,
            in2 => \N__35238\,
            in3 => \N__36384\,
            lcout => \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.periodCounter_RNIV91B_14_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36618\,
            in2 => \_gnd_net_\,
            in3 => \N__36596\,
            lcout => OPEN,
            ltout => \PWMInstance2.un1_periodCounter12_1_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.periodCounter_RNI3BPO_10_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__36576\,
            in1 => \N__36558\,
            in2 => \N__36537\,
            in3 => \N__36219\,
            lcout => \PWMInstance2.un1_periodCounter12_1_0_a2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_4_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36501\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38647\,
            ce => \N__35865\,
            sr => \N__35796\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_5_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36345\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38647\,
            ce => \N__35865\,
            sr => \N__35796\
        );

    \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36218\,
            in1 => \N__35871\,
            in2 => \N__36201\,
            in3 => \N__36021\,
            lcout => \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_10_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36150\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38647\,
            ce => \N__35865\,
            sr => \N__35796\
        );

    \PWMInstance2.PWMPulseWidthCount_esr_11_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36013\,
            lcout => \PWMInstance2.PWMPulseWidthCountZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38647\,
            ce => \N__35865\,
            sr => \N__35796\
        );

    \PWM2_obufLegalizeSB_DFF_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM2_obufLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36916\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM3_obufLegalizeSB_DFF_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM3_obufLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36916\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \MISO_obufLegalizeSB_DFF_LC_20_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \MISO_obufLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_2_5_LC_20_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__36873\,
            in1 => \N__38158\,
            in2 => \N__36831\,
            in3 => \N__36795\,
            lcout => \OutReg_ess_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_1_5_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__36783\,
            in1 => \N__37759\,
            in2 => \N__36750\,
            in3 => \N__36711\,
            lcout => OPEN,
            ltout => \OutReg_ess_RNO_1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_0_5_LC_20_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37565\,
            in2 => \N__36696\,
            in3 => \N__36693\,
            lcout => \OutReg_ess_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_5_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__38901\,
            in1 => \N__36687\,
            in2 => \N__36681\,
            in3 => \N__37387\,
            lcout => \OutRegZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38714\,
            ce => \N__37243\,
            sr => \N__37137\
        );

    \dataOut_RNO_0_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110011"
        )
    port map (
            in0 => \N__39053\,
            in1 => \N__38864\,
            in2 => \N__39090\,
            in3 => \N__37344\,
            lcout => OPEN,
            ltout => \dataOut_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dataOut_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001010"
        )
    port map (
            in0 => \N__36654\,
            in1 => \N__36629\,
            in2 => \N__36642\,
            in3 => \N__39056\,
            lcout => \MISO_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SSELr_0_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37863\,
            lcout => \SSELrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_RNI8CK3_0_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__37810\,
            in1 => \N__38760\,
            in2 => \_gnd_net_\,
            in3 => \N__38798\,
            lcout => un1_bit_count_1_c1,
            ltout => \un1_bit_count_1_c1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_2_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__39054\,
            in1 => \N__37887\,
            in2 => \N__37845\,
            in3 => \N__37962\,
            lcout => \bit_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_ess_RNO_0_15_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37564\,
            in1 => \N__37842\,
            in2 => \_gnd_net_\,
            in3 => \N__37830\,
            lcout => \OutReg_ess_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_0_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100110"
        )
    port map (
            in0 => \N__37811\,
            in1 => \N__38761\,
            in2 => \N__38805\,
            in3 => \N__39055\,
            lcout => \bit_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_1_8_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__37794\,
            in1 => \N__37760\,
            in2 => \N__37617\,
            in3 => \N__37578\,
            lcout => OPEN,
            ltout => \OutReg_esr_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_RNO_0_8_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37569\,
            in1 => \_gnd_net_\,
            in2 => \N__37410\,
            in3 => \N__38001\,
            lcout => OPEN,
            ltout => \OutReg_esr_RNO_0Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutReg_esr_8_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__37407\,
            in1 => \N__38865\,
            in2 => \N__37398\,
            in3 => \N__37381\,
            lcout => \OutRegZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38701\,
            ce => \N__37240\,
            sr => \N__37134\
        );

    \OutReg_esr_RNO_2_8_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__37017\,
            in1 => \N__36980\,
            in2 => \N__38166\,
            in3 => \N__38013\,
            lcout => \OutReg_esr_RNO_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SSELr_1_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37995\,
            lcout => \SSELrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SSELr_2_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39046\,
            lcout => \SSELrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SCKr_0_LC_21_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37971\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \SCKrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38724\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_RNI9MD6_2_LC_21_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__37895\,
            in1 => \N__37960\,
            in2 => \_gnd_net_\,
            in3 => \N__37884\,
            lcout => un1_bit_count_1_c3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SCKr_RNIBA7C_2_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__39047\,
            in1 => \N__38758\,
            in2 => \_gnd_net_\,
            in3 => \N__38796\,
            lcout => \SCKr_RNIBA7CZ0Z_2\,
            ltout => \SCKr_RNIBA7CZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SCKr_RNIMKEO_2_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__38797\,
            in1 => \N__38759\,
            in2 => \N__37926\,
            in3 => \N__39048\,
            lcout => \N_45_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SCKr_1_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37905\,
            lcout => \SCKrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_1_LC_21_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__37896\,
            in1 => \N__39049\,
            in2 => \_gnd_net_\,
            in3 => \N__37885\,
            lcout => \bit_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_4_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__38967\,
            in1 => \N__39036\,
            in2 => \N__38997\,
            in3 => \N__38985\,
            lcout => \bit_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_RNIU615_0_4_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011111"
        )
    port map (
            in0 => \N__38966\,
            in1 => \N__38794\,
            in2 => \N__38763\,
            in3 => \N__38983\,
            lcout => \bit_count_RNIU615_0Z0Z_4\,
            ltout => \bit_count_RNIU615_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SSELr_RNIGO0F_1_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39081\,
            in3 => \N__39034\,
            lcout => \SSELr_RNIGO0FZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_3_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39035\,
            in1 => \N__38993\,
            in2 => \_gnd_net_\,
            in3 => \N__38984\,
            lcout => \bit_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \bit_count_RNIU615_4_LC_21_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__38982\,
            in1 => \N__38965\,
            in2 => \N__38762\,
            in3 => \N__38793\,
            lcout => \un1_OutReg51_4_0_i_o3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SCKr_2_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38795\,
            lcout => \SCKrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38709\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
